// This is the unpowered netlist.
module lifo (clk,
    empty,
    error,
    full,
    pop,
    push,
    rst,
    data_in,
    data_out);
 input clk;
 output empty;
 output error;
 output full;
 input pop;
 input push;
 input rst;
 input [7:0] data_in;
 output [7:0] data_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \stack[0][0] ;
 wire \stack[0][1] ;
 wire \stack[0][2] ;
 wire \stack[0][3] ;
 wire \stack[0][4] ;
 wire \stack[0][5] ;
 wire \stack[0][6] ;
 wire \stack[0][7] ;
 wire \stack[10][0] ;
 wire \stack[10][1] ;
 wire \stack[10][2] ;
 wire \stack[10][3] ;
 wire \stack[10][4] ;
 wire \stack[10][5] ;
 wire \stack[10][6] ;
 wire \stack[10][7] ;
 wire \stack[11][0] ;
 wire \stack[11][1] ;
 wire \stack[11][2] ;
 wire \stack[11][3] ;
 wire \stack[11][4] ;
 wire \stack[11][5] ;
 wire \stack[11][6] ;
 wire \stack[11][7] ;
 wire \stack[12][0] ;
 wire \stack[12][1] ;
 wire \stack[12][2] ;
 wire \stack[12][3] ;
 wire \stack[12][4] ;
 wire \stack[12][5] ;
 wire \stack[12][6] ;
 wire \stack[12][7] ;
 wire \stack[13][0] ;
 wire \stack[13][1] ;
 wire \stack[13][2] ;
 wire \stack[13][3] ;
 wire \stack[13][4] ;
 wire \stack[13][5] ;
 wire \stack[13][6] ;
 wire \stack[13][7] ;
 wire \stack[14][0] ;
 wire \stack[14][1] ;
 wire \stack[14][2] ;
 wire \stack[14][3] ;
 wire \stack[14][4] ;
 wire \stack[14][5] ;
 wire \stack[14][6] ;
 wire \stack[14][7] ;
 wire \stack[15][0] ;
 wire \stack[15][1] ;
 wire \stack[15][2] ;
 wire \stack[15][3] ;
 wire \stack[15][4] ;
 wire \stack[15][5] ;
 wire \stack[15][6] ;
 wire \stack[15][7] ;
 wire \stack[1][0] ;
 wire \stack[1][1] ;
 wire \stack[1][2] ;
 wire \stack[1][3] ;
 wire \stack[1][4] ;
 wire \stack[1][5] ;
 wire \stack[1][6] ;
 wire \stack[1][7] ;
 wire \stack[2][0] ;
 wire \stack[2][1] ;
 wire \stack[2][2] ;
 wire \stack[2][3] ;
 wire \stack[2][4] ;
 wire \stack[2][5] ;
 wire \stack[2][6] ;
 wire \stack[2][7] ;
 wire \stack[3][0] ;
 wire \stack[3][1] ;
 wire \stack[3][2] ;
 wire \stack[3][3] ;
 wire \stack[3][4] ;
 wire \stack[3][5] ;
 wire \stack[3][6] ;
 wire \stack[3][7] ;
 wire \stack[4][0] ;
 wire \stack[4][1] ;
 wire \stack[4][2] ;
 wire \stack[4][3] ;
 wire \stack[4][4] ;
 wire \stack[4][5] ;
 wire \stack[4][6] ;
 wire \stack[4][7] ;
 wire \stack[5][0] ;
 wire \stack[5][1] ;
 wire \stack[5][2] ;
 wire \stack[5][3] ;
 wire \stack[5][4] ;
 wire \stack[5][5] ;
 wire \stack[5][6] ;
 wire \stack[5][7] ;
 wire \stack[6][0] ;
 wire \stack[6][1] ;
 wire \stack[6][2] ;
 wire \stack[6][3] ;
 wire \stack[6][4] ;
 wire \stack[6][5] ;
 wire \stack[6][6] ;
 wire \stack[6][7] ;
 wire \stack[7][0] ;
 wire \stack[7][1] ;
 wire \stack[7][2] ;
 wire \stack[7][3] ;
 wire \stack[7][4] ;
 wire \stack[7][5] ;
 wire \stack[7][6] ;
 wire \stack[7][7] ;
 wire \stack[8][0] ;
 wire \stack[8][1] ;
 wire \stack[8][2] ;
 wire \stack[8][3] ;
 wire \stack[8][4] ;
 wire \stack[8][5] ;
 wire \stack[8][6] ;
 wire \stack[8][7] ;
 wire \stack[9][0] ;
 wire \stack[9][1] ;
 wire \stack[9][2] ;
 wire \stack[9][3] ;
 wire \stack[9][4] ;
 wire \stack[9][5] ;
 wire \stack[9][6] ;
 wire \stack[9][7] ;
 wire \top[0] ;
 wire \top[1] ;
 wire \top[2] ;
 wire \top[3] ;
 wire \top[4] ;

 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__or4_4 _0480_ (.A(\top[3] ),
    .B(\top[2] ),
    .C(\top[1] ),
    .D(\top[0] ),
    .X(_0155_));
 sky130_fd_sc_hd__o21ai_4 _0481_ (.A1(\top[4] ),
    .A2(_0155_),
    .B1(net9),
    .Y(_0156_));
 sky130_fd_sc_hd__buf_2 _0482_ (.A(\top[3] ),
    .X(_0157_));
 sky130_fd_sc_hd__nor4_1 _0483_ (.A(_0157_),
    .B(\top[2] ),
    .C(\top[1] ),
    .D(\top[0] ),
    .Y(_0158_));
 sky130_fd_sc_hd__clkbuf_4 _0484_ (.A(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_4 _0485_ (.A(\top[0] ),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_2 _0486_ (.A(\top[2] ),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_2 _0487_ (.A(\top[1] ),
    .X(_0162_));
 sky130_fd_sc_hd__or3b_2 _0488_ (.A(_0157_),
    .B(_0161_),
    .C_N(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_4 _0489_ (.A(_0160_),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__buf_2 _0490_ (.A(\top[0] ),
    .X(_0165_));
 sky130_fd_sc_hd__and4b_1 _0491_ (.A_N(_0157_),
    .B(_0161_),
    .C(_0162_),
    .D(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _0492_ (.A(_0166_),
    .X(_0167_));
 sky130_fd_sc_hd__buf_2 _0493_ (.A(_0157_),
    .X(_0168_));
 sky130_fd_sc_hd__and4_1 _0494_ (.A(_0168_),
    .B(_0161_),
    .C(_0162_),
    .D(_0165_),
    .X(_0169_));
 sky130_fd_sc_hd__clkbuf_4 _0495_ (.A(_0169_),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _0496_ (.A1(\stack[6][7] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][7] ),
    .X(_0171_));
 sky130_fd_sc_hd__a221o_1 _0497_ (.A1(\stack[15][7] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][7] ),
    .C1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_4 _0498_ (.A(_0162_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_2 _0499_ (.A(_0161_),
    .X(_0174_));
 sky130_fd_sc_hd__and4bb_4 _0500_ (.A_N(_0168_),
    .B_N(_0173_),
    .C(_0160_),
    .D(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(_0165_),
    .Y(_0176_));
 sky130_fd_sc_hd__nor2_4 _0502_ (.A(_0176_),
    .B(_0163_),
    .Y(_0177_));
 sky130_fd_sc_hd__and4b_1 _0503_ (.A_N(_0161_),
    .B(_0162_),
    .C(_0165_),
    .D(_0157_),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_4 _0504_ (.A(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__and4bb_4 _0505_ (.A_N(_0173_),
    .B_N(_0160_),
    .C(_0168_),
    .D(_0174_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _0506_ (.A1(\stack[10][7] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][7] ),
    .X(_0181_));
 sky130_fd_sc_hd__a221o_1 _0507_ (.A1(\stack[4][7] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][7] ),
    .C1(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__nor4b_1 _0508_ (.A(_0161_),
    .B(_0173_),
    .C(_0165_),
    .D_N(_0157_),
    .Y(_0183_));
 sky130_fd_sc_hd__and4b_1 _0509_ (.A_N(_0162_),
    .B(_0165_),
    .C(_0157_),
    .D(_0161_),
    .X(_0184_));
 sky130_fd_sc_hd__clkbuf_4 _0510_ (.A(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _0511_ (.A1(\stack[7][7] ),
    .A2(net28),
    .B1(_0185_),
    .B2(\stack[12][7] ),
    .X(_0186_));
 sky130_fd_sc_hd__and4bb_4 _0512_ (.A_N(_0161_),
    .B_N(_0173_),
    .C(_0165_),
    .D(_0157_),
    .X(_0187_));
 sky130_fd_sc_hd__and4bb_4 _0513_ (.A_N(_0174_),
    .B_N(_0165_),
    .C(_0162_),
    .D(_0157_),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _0514_ (.A1(\stack[8][7] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][7] ),
    .X(_0189_));
 sky130_fd_sc_hd__and4bb_4 _0515_ (.A_N(_0168_),
    .B_N(_0160_),
    .C(_0162_),
    .D(_0161_),
    .X(_0190_));
 sky130_fd_sc_hd__nor4b_2 _0516_ (.A(_0168_),
    .B(_0174_),
    .C(_0173_),
    .D_N(_0160_),
    .Y(_0191_));
 sky130_fd_sc_hd__a21o_1 _0517_ (.A1(\stack[5][7] ),
    .A2(_0190_),
    .B1(net26),
    .X(_0192_));
 sky130_fd_sc_hd__nor4b_2 _0518_ (.A(_0168_),
    .B(_0173_),
    .C(_0160_),
    .D_N(_0174_),
    .Y(_0193_));
 sky130_fd_sc_hd__and4b_1 _0519_ (.A_N(_0165_),
    .B(_0162_),
    .C(_0161_),
    .D(_0157_),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_4 _0520_ (.A(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _0521_ (.A1(\stack[3][7] ),
    .A2(net24),
    .B1(_0195_),
    .B2(\stack[13][7] ),
    .X(_0196_));
 sky130_fd_sc_hd__or4_1 _0522_ (.A(_0186_),
    .B(_0189_),
    .C(_0192_),
    .D(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__or3_1 _0523_ (.A(_0172_),
    .B(_0182_),
    .C(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__or4_4 _0524_ (.A(_0168_),
    .B(_0174_),
    .C(_0173_),
    .D(_0176_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(net9),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_2 _0526_ (.A(\top[4] ),
    .B(_0155_),
    .Y(net20));
 sky130_fd_sc_hd__nor2_4 _0527_ (.A(_0200_),
    .B(net20),
    .Y(_0201_));
 sky130_fd_sc_hd__o21a_1 _0528_ (.A1(net148),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _0529_ (.A1(net159),
    .A2(_0156_),
    .B1(_0198_),
    .B2(_0202_),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _0530_ (.A1(\stack[6][6] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][6] ),
    .X(_0203_));
 sky130_fd_sc_hd__a221o_1 _0531_ (.A1(\stack[15][6] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][6] ),
    .C1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _0532_ (.A1(\stack[10][6] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][6] ),
    .X(_0205_));
 sky130_fd_sc_hd__a221o_1 _0533_ (.A1(\stack[4][6] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][6] ),
    .C1(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _0534_ (.A1(\stack[7][6] ),
    .A2(net28),
    .B1(_0185_),
    .B2(\stack[12][6] ),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_1 _0535_ (.A1(\stack[8][6] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][6] ),
    .X(_0208_));
 sky130_fd_sc_hd__a21o_1 _0536_ (.A1(\stack[5][6] ),
    .A2(_0190_),
    .B1(net26),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _0537_ (.A1(\stack[3][6] ),
    .A2(net24),
    .B1(_0195_),
    .B2(\stack[13][6] ),
    .X(_0210_));
 sky130_fd_sc_hd__or4_1 _0538_ (.A(_0207_),
    .B(_0208_),
    .C(_0209_),
    .D(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__or3_1 _0539_ (.A(_0204_),
    .B(_0206_),
    .C(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__o21a_1 _0540_ (.A1(\stack[0][6] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _0541_ (.A1(net34),
    .A2(_0156_),
    .B1(_0212_),
    .B2(_0213_),
    .X(_0033_));
 sky130_fd_sc_hd__a22o_1 _0542_ (.A1(\stack[6][5] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][5] ),
    .X(_0214_));
 sky130_fd_sc_hd__a221o_1 _0543_ (.A1(\stack[15][5] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][5] ),
    .C1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _0544_ (.A1(\stack[10][5] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][5] ),
    .X(_0216_));
 sky130_fd_sc_hd__a221o_1 _0545_ (.A1(\stack[4][5] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][5] ),
    .C1(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _0546_ (.A1(\stack[7][5] ),
    .A2(net27),
    .B1(_0185_),
    .B2(\stack[12][5] ),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _0547_ (.A1(\stack[8][5] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][5] ),
    .X(_0219_));
 sky130_fd_sc_hd__a21o_1 _0548_ (.A1(\stack[5][5] ),
    .A2(_0190_),
    .B1(net25),
    .X(_0220_));
 sky130_fd_sc_hd__a22o_1 _0549_ (.A1(\stack[3][5] ),
    .A2(net23),
    .B1(_0195_),
    .B2(\stack[13][5] ),
    .X(_0221_));
 sky130_fd_sc_hd__or4_1 _0550_ (.A(_0218_),
    .B(_0219_),
    .C(_0220_),
    .D(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__or3_1 _0551_ (.A(_0215_),
    .B(_0217_),
    .C(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__o21a_1 _0552_ (.A1(\stack[0][5] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0224_));
 sky130_fd_sc_hd__a22o_1 _0553_ (.A1(net42),
    .A2(_0156_),
    .B1(_0223_),
    .B2(_0224_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _0554_ (.A1(\stack[6][4] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][4] ),
    .X(_0225_));
 sky130_fd_sc_hd__a221o_1 _0555_ (.A1(\stack[15][4] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][4] ),
    .C1(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _0556_ (.A1(\stack[10][4] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][4] ),
    .X(_0227_));
 sky130_fd_sc_hd__a221o_1 _0557_ (.A1(\stack[4][4] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][4] ),
    .C1(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _0558_ (.A1(\stack[7][4] ),
    .A2(net28),
    .B1(_0185_),
    .B2(\stack[12][4] ),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _0559_ (.A1(\stack[8][4] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][4] ),
    .X(_0230_));
 sky130_fd_sc_hd__a21o_1 _0560_ (.A1(\stack[5][4] ),
    .A2(_0190_),
    .B1(net26),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _0561_ (.A1(\stack[3][4] ),
    .A2(net24),
    .B1(_0195_),
    .B2(\stack[13][4] ),
    .X(_0232_));
 sky130_fd_sc_hd__or4_2 _0562_ (.A(_0229_),
    .B(_0230_),
    .C(_0231_),
    .D(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__or3_1 _0563_ (.A(_0226_),
    .B(_0228_),
    .C(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__o21a_1 _0564_ (.A1(\stack[0][4] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _0565_ (.A1(net32),
    .A2(_0156_),
    .B1(_0234_),
    .B2(_0235_),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _0566_ (.A1(\stack[6][3] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][3] ),
    .X(_0236_));
 sky130_fd_sc_hd__a221o_1 _0567_ (.A1(\stack[15][3] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][3] ),
    .C1(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_1 _0568_ (.A1(\stack[10][3] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][3] ),
    .X(_0238_));
 sky130_fd_sc_hd__a221o_1 _0569_ (.A1(\stack[4][3] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][3] ),
    .C1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _0570_ (.A1(\stack[7][3] ),
    .A2(net27),
    .B1(_0185_),
    .B2(\stack[12][3] ),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _0571_ (.A1(\stack[8][3] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][3] ),
    .X(_0241_));
 sky130_fd_sc_hd__a21o_1 _0572_ (.A1(\stack[5][3] ),
    .A2(_0190_),
    .B1(net25),
    .X(_0242_));
 sky130_fd_sc_hd__a22o_1 _0573_ (.A1(\stack[3][3] ),
    .A2(net23),
    .B1(_0195_),
    .B2(\stack[13][3] ),
    .X(_0243_));
 sky130_fd_sc_hd__or4_1 _0574_ (.A(_0240_),
    .B(_0241_),
    .C(_0242_),
    .D(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__or3_1 _0575_ (.A(_0237_),
    .B(_0239_),
    .C(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__o21a_1 _0576_ (.A1(\stack[0][3] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _0577_ (.A1(net38),
    .A2(_0156_),
    .B1(_0245_),
    .B2(_0246_),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _0578_ (.A1(\stack[6][2] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][2] ),
    .X(_0247_));
 sky130_fd_sc_hd__a221o_1 _0579_ (.A1(\stack[15][2] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][2] ),
    .C1(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _0580_ (.A1(\stack[10][2] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][2] ),
    .X(_0249_));
 sky130_fd_sc_hd__a221o_1 _0581_ (.A1(\stack[4][2] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][2] ),
    .C1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _0582_ (.A1(\stack[7][2] ),
    .A2(net27),
    .B1(_0185_),
    .B2(\stack[12][2] ),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _0583_ (.A1(\stack[8][2] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][2] ),
    .X(_0252_));
 sky130_fd_sc_hd__a21o_1 _0584_ (.A1(\stack[5][2] ),
    .A2(_0190_),
    .B1(net25),
    .X(_0253_));
 sky130_fd_sc_hd__a22o_1 _0585_ (.A1(\stack[3][2] ),
    .A2(net23),
    .B1(_0195_),
    .B2(\stack[13][2] ),
    .X(_0254_));
 sky130_fd_sc_hd__or4_1 _0586_ (.A(_0251_),
    .B(_0252_),
    .C(_0253_),
    .D(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__or3_1 _0587_ (.A(_0248_),
    .B(_0250_),
    .C(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__o21a_1 _0588_ (.A1(\stack[0][2] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _0589_ (.A1(net36),
    .A2(_0156_),
    .B1(_0256_),
    .B2(_0257_),
    .X(_0029_));
 sky130_fd_sc_hd__a22o_1 _0590_ (.A1(\stack[6][1] ),
    .A2(_0167_),
    .B1(_0170_),
    .B2(\stack[14][1] ),
    .X(_0258_));
 sky130_fd_sc_hd__a221o_1 _0591_ (.A1(\stack[15][1] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][1] ),
    .C1(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _0592_ (.A1(\stack[10][1] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][1] ),
    .X(_0260_));
 sky130_fd_sc_hd__a221o_1 _0593_ (.A1(\stack[4][1] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][1] ),
    .C1(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _0594_ (.A1(\stack[7][1] ),
    .A2(net27),
    .B1(_0185_),
    .B2(\stack[12][1] ),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _0595_ (.A1(\stack[8][1] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][1] ),
    .X(_0263_));
 sky130_fd_sc_hd__a21o_1 _0596_ (.A1(\stack[5][1] ),
    .A2(_0190_),
    .B1(net25),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _0597_ (.A1(\stack[3][1] ),
    .A2(net23),
    .B1(_0195_),
    .B2(\stack[13][1] ),
    .X(_0265_));
 sky130_fd_sc_hd__or4_1 _0598_ (.A(_0262_),
    .B(_0263_),
    .C(_0264_),
    .D(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__or3_1 _0599_ (.A(_0259_),
    .B(_0261_),
    .C(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__o21a_1 _0600_ (.A1(\stack[0][1] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _0601_ (.A1(net112),
    .A2(_0156_),
    .B1(_0267_),
    .B2(_0268_),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_1 _0602_ (.A1(\stack[6][0] ),
    .A2(_0167_),
    .B1(_0169_),
    .B2(\stack[14][0] ),
    .X(_0269_));
 sky130_fd_sc_hd__a221o_1 _0603_ (.A1(\stack[15][0] ),
    .A2(_0159_),
    .B1(_0164_),
    .B2(\stack[1][0] ),
    .C1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _0604_ (.A1(\stack[10][0] ),
    .A2(_0179_),
    .B1(_0180_),
    .B2(\stack[11][0] ),
    .X(_0271_));
 sky130_fd_sc_hd__a221o_1 _0605_ (.A1(\stack[4][0] ),
    .A2(_0175_),
    .B1(_0177_),
    .B2(\stack[2][0] ),
    .C1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _0606_ (.A1(\stack[7][0] ),
    .A2(net27),
    .B1(_0185_),
    .B2(\stack[12][0] ),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _0607_ (.A1(\stack[8][0] ),
    .A2(_0187_),
    .B1(_0188_),
    .B2(\stack[9][0] ),
    .X(_0274_));
 sky130_fd_sc_hd__a21o_1 _0608_ (.A1(\stack[5][0] ),
    .A2(_0190_),
    .B1(net26),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _0609_ (.A1(\stack[3][0] ),
    .A2(net23),
    .B1(_0195_),
    .B2(\stack[13][0] ),
    .X(_0276_));
 sky130_fd_sc_hd__or4_1 _0610_ (.A(_0273_),
    .B(_0274_),
    .C(_0275_),
    .D(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__or3_1 _0611_ (.A(_0270_),
    .B(_0272_),
    .C(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__o21a_1 _0612_ (.A1(\stack[0][0] ),
    .A2(_0199_),
    .B1(_0201_),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_1 _0613_ (.A1(net30),
    .A2(_0156_),
    .B1(_0278_),
    .B2(_0279_),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _0614_ (.A(_0200_),
    .B(net10),
    .C(_0170_),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_1 _0615_ (.A1(net9),
    .A2(_0159_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__mux2_1 _0616_ (.A0(_0280_),
    .A1(_0281_),
    .S(\top[4] ),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_1 _0617_ (.A(_0282_),
    .X(_0026_));
 sky130_fd_sc_hd__or2_1 _0618_ (.A(_0162_),
    .B(_0165_),
    .X(_0283_));
 sky130_fd_sc_hd__or2_1 _0619_ (.A(_0174_),
    .B(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _0620_ (.A(\top[4] ),
    .B(_0159_),
    .X(_0285_));
 sky130_fd_sc_hd__buf_1 _0621_ (.A(_0285_),
    .X(net22));
 sky130_fd_sc_hd__a21o_1 _0622_ (.A1(_0168_),
    .A2(_0284_),
    .B1(net22),
    .X(_0286_));
 sky130_fd_sc_hd__a31o_1 _0623_ (.A1(_0174_),
    .A2(_0173_),
    .A3(_0160_),
    .B1(_0168_),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_1 _0624_ (.A(net9),
    .B(_0170_),
    .Y(_0288_));
 sky130_fd_sc_hd__a22o_1 _0625_ (.A1(net9),
    .A2(_0286_),
    .B1(_0287_),
    .B2(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__inv_2 _0626_ (.A(net10),
    .Y(_0290_));
 sky130_fd_sc_hd__and3_1 _0627_ (.A(net9),
    .B(net10),
    .C(_0155_),
    .X(_0291_));
 sky130_fd_sc_hd__buf_2 _0628_ (.A(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__a21oi_2 _0629_ (.A1(_0290_),
    .A2(_0156_),
    .B1(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__mux2_1 _0630_ (.A0(_0168_),
    .A1(_0289_),
    .S(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _0631_ (.A(_0294_),
    .X(_0025_));
 sky130_fd_sc_hd__nand2_1 _0632_ (.A(_0173_),
    .B(_0160_),
    .Y(_0295_));
 sky130_fd_sc_hd__xor2_1 _0633_ (.A(_0174_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__a21oi_1 _0634_ (.A1(_0283_),
    .A2(_0295_),
    .B1(_0156_),
    .Y(_0297_));
 sky130_fd_sc_hd__xnor2_1 _0635_ (.A(_0296_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_1 _0636_ (.A0(_0174_),
    .A1(_0298_),
    .S(_0293_),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_1 _0637_ (.A(_0299_),
    .X(_0024_));
 sky130_fd_sc_hd__a31o_1 _0638_ (.A1(_0200_),
    .A2(_0283_),
    .A3(_0295_),
    .B1(_0297_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _0639_ (.A0(_0173_),
    .A1(_0300_),
    .S(_0293_),
    .X(_0301_));
 sky130_fd_sc_hd__clkbuf_1 _0640_ (.A(_0301_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _0641_ (.A(_0200_),
    .B(net10),
    .C(net22),
    .X(_0302_));
 sky130_fd_sc_hd__nor2_1 _0642_ (.A(_0160_),
    .B(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hd__mux2_1 _0643_ (.A0(_0160_),
    .A1(_0303_),
    .S(_0293_),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(_0304_),
    .X(_0022_));
 sky130_fd_sc_hd__a31o_1 _0645_ (.A1(net9),
    .A2(_0290_),
    .A3(net20),
    .B1(_0302_),
    .X(_0479_));
 sky130_fd_sc_hd__clkbuf_4 _0646_ (.A(net1),
    .X(_0305_));
 sky130_fd_sc_hd__inv_2 _0647_ (.A(net11),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_4 _0648_ (.A(_0000_),
    .B(_0280_),
    .Y(_0306_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(_0305_),
    .A1(net133),
    .S(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0307_),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_4 _0651_ (.A(net2),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _0652_ (.A0(_0308_),
    .A1(net130),
    .S(_0306_),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_1 _0653_ (.A(_0309_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_2 _0654_ (.A(net3),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _0655_ (.A0(_0310_),
    .A1(net168),
    .S(_0306_),
    .X(_0311_));
 sky130_fd_sc_hd__clkbuf_1 _0656_ (.A(_0311_),
    .X(_0016_));
 sky130_fd_sc_hd__buf_2 _0657_ (.A(net4),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _0658_ (.A0(_0312_),
    .A1(net118),
    .S(_0306_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_1 _0659_ (.A(_0313_),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _0660_ (.A(net5),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _0661_ (.A0(_0314_),
    .A1(net161),
    .S(_0306_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_1 _0662_ (.A(_0315_),
    .X(_0018_));
 sky130_fd_sc_hd__buf_2 _0663_ (.A(net6),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _0664_ (.A0(_0316_),
    .A1(net111),
    .S(_0306_),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _0665_ (.A(_0317_),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_4 _0666_ (.A(net7),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(_0318_),
    .A1(net147),
    .S(_0306_),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_1 _0668_ (.A(_0319_),
    .X(_0020_));
 sky130_fd_sc_hd__buf_2 _0669_ (.A(net8),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _0670_ (.A0(_0320_),
    .A1(net152),
    .S(_0306_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _0671_ (.A(_0321_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_8 _0672_ (.A(net11),
    .X(_0322_));
 sky130_fd_sc_hd__inv_2 _0673_ (.A(_0322_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _0674_ (.A(_0322_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _0675_ (.A(_0322_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _0676_ (.A(_0322_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0677_ (.A(_0322_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _0678_ (.A(_0322_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _0679_ (.A(_0322_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _0680_ (.A(_0322_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(_0322_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _0682_ (.A(_0322_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(net11),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _0684_ (.A(net11),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _0685_ (.A(net11),
    .Y(_0013_));
 sky130_fd_sc_hd__nor2_4 _0686_ (.A(_0290_),
    .B(net11),
    .Y(_0323_));
 sky130_fd_sc_hd__clkbuf_8 _0687_ (.A(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__a21o_1 _0688_ (.A1(_0191_),
    .A2(_0292_),
    .B1(net20),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_4 _0689_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__mux2_1 _0690_ (.A0(_0305_),
    .A1(net122),
    .S(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_1 _0691_ (.A(_0327_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0692_ (.A0(_0308_),
    .A1(net135),
    .S(_0326_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_1 _0693_ (.A(_0328_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _0694_ (.A0(_0310_),
    .A1(net103),
    .S(_0326_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _0695_ (.A(_0329_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0696_ (.A0(_0312_),
    .A1(net146),
    .S(_0326_),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_1 _0697_ (.A(_0330_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0698_ (.A0(_0314_),
    .A1(net145),
    .S(_0326_),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_1 _0699_ (.A(_0331_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0700_ (.A0(_0316_),
    .A1(net106),
    .S(_0326_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _0701_ (.A(_0332_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _0702_ (.A0(_0318_),
    .A1(net86),
    .S(_0326_),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _0703_ (.A(_0333_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0704_ (.A0(_0320_),
    .A1(net148),
    .S(_0326_),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_1 _0705_ (.A(_0334_),
    .X(_0042_));
 sky130_fd_sc_hd__or3_2 _0706_ (.A(_0200_),
    .B(_0290_),
    .C(net29),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _0707_ (.A0(_0164_),
    .A1(net25),
    .S(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _0708_ (.A(_0324_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__mux2_1 _0709_ (.A0(_0305_),
    .A1(net109),
    .S(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_1 _0710_ (.A(_0338_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0711_ (.A0(_0308_),
    .A1(net172),
    .S(_0337_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0339_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _0713_ (.A0(_0310_),
    .A1(net163),
    .S(_0337_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0340_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0715_ (.A0(_0312_),
    .A1(net164),
    .S(_0337_),
    .X(_0341_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0341_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0717_ (.A0(_0314_),
    .A1(net165),
    .S(_0337_),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _0718_ (.A(_0342_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0719_ (.A0(_0316_),
    .A1(net156),
    .S(_0337_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _0720_ (.A(_0343_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0721_ (.A0(_0318_),
    .A1(net171),
    .S(_0337_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0344_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0723_ (.A0(_0320_),
    .A1(net170),
    .S(_0337_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _0724_ (.A(_0345_),
    .X(_0050_));
 sky130_fd_sc_hd__buf_4 _0725_ (.A(_0335_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _0726_ (.A(_0164_),
    .B(_0292_),
    .X(_0347_));
 sky130_fd_sc_hd__o211a_4 _0727_ (.A1(_0177_),
    .A2(_0346_),
    .B1(_0324_),
    .C1(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _0728_ (.A0(net169),
    .A1(_0305_),
    .S(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _0729_ (.A(_0349_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0730_ (.A0(net119),
    .A1(_0308_),
    .S(_0348_),
    .X(_0350_));
 sky130_fd_sc_hd__clkbuf_1 _0731_ (.A(_0350_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _0732_ (.A0(net87),
    .A1(_0310_),
    .S(_0348_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _0733_ (.A(_0351_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(net104),
    .A1(_0312_),
    .S(_0348_),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_1 _0735_ (.A(_0352_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0736_ (.A0(net95),
    .A1(_0314_),
    .S(_0348_),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_1 _0737_ (.A(_0353_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0738_ (.A0(net107),
    .A1(_0316_),
    .S(_0348_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _0739_ (.A(_0354_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _0740_ (.A0(net129),
    .A1(_0318_),
    .S(_0348_),
    .X(_0355_));
 sky130_fd_sc_hd__clkbuf_1 _0741_ (.A(_0355_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0742_ (.A0(net97),
    .A1(_0320_),
    .S(_0348_),
    .X(_0356_));
 sky130_fd_sc_hd__clkbuf_1 _0743_ (.A(_0356_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0744_ (.A0(_0193_),
    .A1(_0177_),
    .S(_0335_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_4 _0745_ (.A(_0324_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__mux2_1 _0746_ (.A0(_0305_),
    .A1(net157),
    .S(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _0747_ (.A(_0359_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(_0308_),
    .A1(net151),
    .S(_0358_),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _0749_ (.A(_0360_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(_0310_),
    .A1(net120),
    .S(_0358_),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _0751_ (.A(_0361_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0752_ (.A0(_0312_),
    .A1(net150),
    .S(_0358_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _0753_ (.A(_0362_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0754_ (.A0(_0314_),
    .A1(net132),
    .S(_0358_),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _0755_ (.A(_0363_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0756_ (.A0(_0316_),
    .A1(net154),
    .S(_0358_),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _0757_ (.A(_0364_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _0758_ (.A0(_0318_),
    .A1(net142),
    .S(_0358_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _0759_ (.A(_0365_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0760_ (.A0(_0320_),
    .A1(net96),
    .S(_0358_),
    .X(_0366_));
 sky130_fd_sc_hd__clkbuf_1 _0761_ (.A(_0366_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _0762_ (.A(_0193_),
    .B(_0292_),
    .X(_0367_));
 sky130_fd_sc_hd__o211a_4 _0763_ (.A1(_0175_),
    .A2(_0346_),
    .B1(_0324_),
    .C1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _0764_ (.A0(net72),
    .A1(_0305_),
    .S(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _0765_ (.A(_0369_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0766_ (.A0(net57),
    .A1(_0308_),
    .S(_0368_),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _0767_ (.A(_0370_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _0768_ (.A0(net46),
    .A1(_0310_),
    .S(_0368_),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _0769_ (.A(_0371_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0770_ (.A0(net115),
    .A1(_0312_),
    .S(_0368_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _0771_ (.A(_0372_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0772_ (.A0(net166),
    .A1(_0314_),
    .S(_0368_),
    .X(_0373_));
 sky130_fd_sc_hd__clkbuf_1 _0773_ (.A(_0373_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0774_ (.A0(net62),
    .A1(_0316_),
    .S(_0368_),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_1 _0775_ (.A(_0374_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _0776_ (.A0(net53),
    .A1(_0318_),
    .S(_0368_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _0777_ (.A(_0375_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0778_ (.A0(net117),
    .A1(_0320_),
    .S(_0368_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_1 _0779_ (.A(_0376_),
    .X(_0074_));
 sky130_fd_sc_hd__or2_1 _0780_ (.A(_0175_),
    .B(_0292_),
    .X(_0377_));
 sky130_fd_sc_hd__o211a_4 _0781_ (.A1(_0190_),
    .A2(_0346_),
    .B1(_0324_),
    .C1(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(net78),
    .A1(_0305_),
    .S(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _0783_ (.A(_0379_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0784_ (.A0(net69),
    .A1(_0308_),
    .S(_0378_),
    .X(_0380_));
 sky130_fd_sc_hd__clkbuf_1 _0785_ (.A(_0380_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _0786_ (.A0(net71),
    .A1(_0310_),
    .S(_0378_),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_1 _0787_ (.A(_0381_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0788_ (.A0(net67),
    .A1(_0312_),
    .S(_0378_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _0789_ (.A(_0382_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0790_ (.A0(net91),
    .A1(_0314_),
    .S(_0378_),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_1 _0791_ (.A(_0383_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0792_ (.A0(net66),
    .A1(_0316_),
    .S(_0378_),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_1 _0793_ (.A(_0384_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0794_ (.A0(net61),
    .A1(_0318_),
    .S(_0378_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_1 _0795_ (.A(_0385_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0796_ (.A0(net85),
    .A1(_0320_),
    .S(_0378_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _0797_ (.A(_0386_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _0798_ (.A0(_0167_),
    .A1(_0190_),
    .S(_0335_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_4 _0799_ (.A(_0324_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__mux2_1 _0800_ (.A0(_0305_),
    .A1(net138),
    .S(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _0801_ (.A(_0389_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0802_ (.A0(_0308_),
    .A1(net123),
    .S(_0388_),
    .X(_0390_));
 sky130_fd_sc_hd__clkbuf_1 _0803_ (.A(_0390_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _0804_ (.A0(_0310_),
    .A1(net136),
    .S(_0388_),
    .X(_0391_));
 sky130_fd_sc_hd__clkbuf_1 _0805_ (.A(_0391_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _0806_ (.A0(_0312_),
    .A1(net110),
    .S(_0388_),
    .X(_0392_));
 sky130_fd_sc_hd__clkbuf_1 _0807_ (.A(_0392_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _0808_ (.A0(_0314_),
    .A1(net167),
    .S(_0388_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _0809_ (.A(_0393_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _0810_ (.A0(_0316_),
    .A1(net101),
    .S(_0388_),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _0811_ (.A(_0394_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _0812_ (.A0(_0318_),
    .A1(net131),
    .S(_0388_),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _0813_ (.A(_0395_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _0814_ (.A0(_0320_),
    .A1(net162),
    .S(_0388_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _0815_ (.A(_0396_),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_1 _0816_ (.A1(net9),
    .A2(_0155_),
    .B1(_0167_),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _0817_ (.A(net9),
    .B(_0284_),
    .Y(_0398_));
 sky130_fd_sc_hd__and3_1 _0818_ (.A(_0323_),
    .B(_0397_),
    .C(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _0819_ (.A(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _0820_ (.A0(net81),
    .A1(_0305_),
    .S(_0400_),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _0821_ (.A(_0401_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _0822_ (.A0(net102),
    .A1(_0308_),
    .S(_0400_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _0823_ (.A(_0402_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _0824_ (.A0(net54),
    .A1(_0310_),
    .S(_0400_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _0825_ (.A(_0403_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _0826_ (.A0(net55),
    .A1(_0312_),
    .S(_0400_),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _0827_ (.A(_0404_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0828_ (.A0(net83),
    .A1(_0314_),
    .S(_0400_),
    .X(_0405_));
 sky130_fd_sc_hd__clkbuf_1 _0829_ (.A(_0405_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _0830_ (.A0(net124),
    .A1(_0316_),
    .S(_0400_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _0831_ (.A(_0406_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _0832_ (.A0(net44),
    .A1(_0318_),
    .S(_0400_),
    .X(_0407_));
 sky130_fd_sc_hd__clkbuf_1 _0833_ (.A(_0407_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _0834_ (.A0(net79),
    .A1(_0320_),
    .S(_0400_),
    .X(_0408_));
 sky130_fd_sc_hd__clkbuf_1 _0835_ (.A(_0408_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _0836_ (.A(_0187_),
    .B(_0346_),
    .X(_0409_));
 sky130_fd_sc_hd__o211a_4 _0837_ (.A1(net173),
    .A2(_0292_),
    .B1(_0324_),
    .C1(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _0838_ (.A0(net52),
    .A1(_0305_),
    .S(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__clkbuf_1 _0839_ (.A(_0411_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _0840_ (.A0(net50),
    .A1(_0308_),
    .S(_0410_),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_1 _0841_ (.A(_0412_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _0842_ (.A0(net92),
    .A1(_0310_),
    .S(_0410_),
    .X(_0413_));
 sky130_fd_sc_hd__clkbuf_1 _0843_ (.A(_0413_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _0844_ (.A0(net51),
    .A1(_0312_),
    .S(_0410_),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _0845_ (.A(_0414_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _0846_ (.A0(net108),
    .A1(_0314_),
    .S(_0410_),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_1 _0847_ (.A(_0415_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _0848_ (.A0(net75),
    .A1(_0316_),
    .S(_0410_),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_1 _0849_ (.A(_0416_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _0850_ (.A0(net74),
    .A1(_0318_),
    .S(_0410_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_1 _0851_ (.A(_0417_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _0852_ (.A0(net73),
    .A1(_0320_),
    .S(_0410_),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_1 _0853_ (.A(_0418_),
    .X(_0106_));
 sky130_fd_sc_hd__or2_1 _0854_ (.A(_0187_),
    .B(_0292_),
    .X(_0419_));
 sky130_fd_sc_hd__o211a_4 _0855_ (.A1(_0188_),
    .A2(_0346_),
    .B1(_0324_),
    .C1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _0856_ (.A0(net100),
    .A1(net1),
    .S(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _0857_ (.A(_0421_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _0858_ (.A0(net40),
    .A1(net2),
    .S(_0420_),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _0859_ (.A(_0422_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0860_ (.A0(net84),
    .A1(net3),
    .S(_0420_),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _0861_ (.A(_0423_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(net58),
    .A1(net4),
    .S(_0420_),
    .X(_0424_));
 sky130_fd_sc_hd__clkbuf_1 _0863_ (.A(_0424_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _0864_ (.A0(net125),
    .A1(net5),
    .S(_0420_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_1 _0865_ (.A(_0425_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _0866_ (.A0(net93),
    .A1(net6),
    .S(_0420_),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_1 _0867_ (.A(_0426_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _0868_ (.A0(net134),
    .A1(net7),
    .S(_0420_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_1 _0869_ (.A(_0427_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _0870_ (.A0(net45),
    .A1(net8),
    .S(_0420_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_1 _0871_ (.A(_0428_),
    .X(_0114_));
 sky130_fd_sc_hd__or2_1 _0872_ (.A(_0188_),
    .B(_0292_),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_4 _0873_ (.A1(_0179_),
    .A2(_0346_),
    .B1(_0324_),
    .C1(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _0874_ (.A0(net139),
    .A1(net1),
    .S(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_1 _0875_ (.A(_0431_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _0876_ (.A0(net59),
    .A1(net2),
    .S(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_1 _0877_ (.A(_0432_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _0878_ (.A0(net65),
    .A1(net3),
    .S(_0430_),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_1 _0879_ (.A(_0433_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(net126),
    .A1(net4),
    .S(_0430_),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_1 _0881_ (.A(_0434_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0882_ (.A0(net94),
    .A1(net5),
    .S(_0430_),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_1 _0883_ (.A(_0435_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(net77),
    .A1(net6),
    .S(_0430_),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_1 _0885_ (.A(_0436_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(net41),
    .A1(net7),
    .S(_0430_),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_1 _0887_ (.A(_0437_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _0888_ (.A0(net105),
    .A1(net8),
    .S(_0430_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_1 _0889_ (.A(_0438_),
    .X(_0122_));
 sky130_fd_sc_hd__or2_1 _0890_ (.A(_0179_),
    .B(_0292_),
    .X(_0439_));
 sky130_fd_sc_hd__o211a_4 _0891_ (.A1(_0180_),
    .A2(_0346_),
    .B1(_0323_),
    .C1(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(net82),
    .A1(net1),
    .S(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_1 _0893_ (.A(_0441_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0894_ (.A0(net149),
    .A1(net2),
    .S(_0440_),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_1 _0895_ (.A(_0442_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(net76),
    .A1(net3),
    .S(_0440_),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_1 _0897_ (.A(_0443_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(net141),
    .A1(net4),
    .S(_0440_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_1 _0899_ (.A(_0444_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _0900_ (.A0(net63),
    .A1(net5),
    .S(_0440_),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_1 _0901_ (.A(_0445_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(net68),
    .A1(net6),
    .S(_0440_),
    .X(_0446_));
 sky130_fd_sc_hd__clkbuf_1 _0903_ (.A(_0446_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(net80),
    .A1(net7),
    .S(_0440_),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_1 _0905_ (.A(_0447_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(net114),
    .A1(net8),
    .S(_0440_),
    .X(_0448_));
 sky130_fd_sc_hd__clkbuf_1 _0907_ (.A(_0448_),
    .X(_0130_));
 sky130_fd_sc_hd__or2_1 _0908_ (.A(_0180_),
    .B(_0292_),
    .X(_0449_));
 sky130_fd_sc_hd__o211a_4 _0909_ (.A1(_0185_),
    .A2(_0346_),
    .B1(_0323_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(net137),
    .A1(net1),
    .S(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_1 _0911_ (.A(_0451_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(net99),
    .A1(net2),
    .S(_0450_),
    .X(_0452_));
 sky130_fd_sc_hd__clkbuf_1 _0913_ (.A(_0452_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(net158),
    .A1(net3),
    .S(_0450_),
    .X(_0453_));
 sky130_fd_sc_hd__clkbuf_1 _0915_ (.A(_0453_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(net155),
    .A1(net4),
    .S(_0450_),
    .X(_0454_));
 sky130_fd_sc_hd__clkbuf_1 _0917_ (.A(_0454_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(net116),
    .A1(net5),
    .S(_0450_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_1 _0919_ (.A(_0455_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0920_ (.A0(net127),
    .A1(net6),
    .S(_0450_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_1 _0921_ (.A(_0456_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(net144),
    .A1(net7),
    .S(_0450_),
    .X(_0457_));
 sky130_fd_sc_hd__clkbuf_1 _0923_ (.A(_0457_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(net70),
    .A1(net8),
    .S(_0450_),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _0925_ (.A(_0458_),
    .X(_0138_));
 sky130_fd_sc_hd__or2_1 _0926_ (.A(_0185_),
    .B(_0291_),
    .X(_0459_));
 sky130_fd_sc_hd__o211a_4 _0927_ (.A1(_0195_),
    .A2(_0346_),
    .B1(_0323_),
    .C1(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net160),
    .A1(net1),
    .S(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _0929_ (.A(_0461_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(net89),
    .A1(net2),
    .S(_0460_),
    .X(_0462_));
 sky130_fd_sc_hd__clkbuf_1 _0931_ (.A(_0462_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net60),
    .A1(net3),
    .S(_0460_),
    .X(_0463_));
 sky130_fd_sc_hd__clkbuf_1 _0933_ (.A(_0463_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net88),
    .A1(net4),
    .S(_0460_),
    .X(_0464_));
 sky130_fd_sc_hd__clkbuf_1 _0935_ (.A(_0464_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _0936_ (.A0(net121),
    .A1(net5),
    .S(_0460_),
    .X(_0465_));
 sky130_fd_sc_hd__clkbuf_1 _0937_ (.A(_0465_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(net153),
    .A1(net6),
    .S(_0460_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_1 _0939_ (.A(_0466_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(net140),
    .A1(net7),
    .S(_0460_),
    .X(_0467_));
 sky130_fd_sc_hd__clkbuf_1 _0941_ (.A(_0467_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _0942_ (.A0(net56),
    .A1(net8),
    .S(_0460_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_1 _0943_ (.A(_0468_),
    .X(_0146_));
 sky130_fd_sc_hd__or2_1 _0944_ (.A(_0195_),
    .B(_0291_),
    .X(_0469_));
 sky130_fd_sc_hd__o211a_4 _0945_ (.A1(_0170_),
    .A2(_0346_),
    .B1(_0323_),
    .C1(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(net48),
    .A1(net1),
    .S(_0470_),
    .X(_0471_));
 sky130_fd_sc_hd__clkbuf_1 _0947_ (.A(_0471_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(net98),
    .A1(net2),
    .S(_0470_),
    .X(_0472_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0472_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net64),
    .A1(net3),
    .S(_0470_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0473_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _0952_ (.A0(net143),
    .A1(net4),
    .S(_0470_),
    .X(_0474_));
 sky130_fd_sc_hd__clkbuf_1 _0953_ (.A(_0474_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net90),
    .A1(net5),
    .S(_0470_),
    .X(_0475_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0475_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net49),
    .A1(net6),
    .S(_0470_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0476_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(net47),
    .A1(net7),
    .S(_0470_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0477_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net128),
    .A1(net8),
    .S(_0470_),
    .X(_0478_));
 sky130_fd_sc_hd__clkbuf_1 _0961_ (.A(_0478_),
    .X(_0154_));
 sky130_fd_sc_hd__dfxtp_1 _0962_ (.CLK(clknet_4_3_0_clk),
    .D(_0014_),
    .Q(\stack[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0963_ (.CLK(clknet_4_1_0_clk),
    .D(_0015_),
    .Q(\stack[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0964_ (.CLK(clknet_4_1_0_clk),
    .D(_0016_),
    .Q(\stack[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0965_ (.CLK(clknet_4_3_0_clk),
    .D(_0017_),
    .Q(\stack[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0966_ (.CLK(clknet_4_5_0_clk),
    .D(_0018_),
    .Q(\stack[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0967_ (.CLK(clknet_4_3_0_clk),
    .D(_0019_),
    .Q(\stack[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0968_ (.CLK(clknet_4_7_0_clk),
    .D(_0020_),
    .Q(\stack[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0969_ (.CLK(clknet_4_5_0_clk),
    .D(_0021_),
    .Q(\stack[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0970_ (.CLK(clknet_4_7_0_clk),
    .D(_0022_),
    .RESET_B(_0000_),
    .Q(\top[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0971_ (.CLK(clknet_4_7_0_clk),
    .D(_0023_),
    .RESET_B(_0001_),
    .Q(\top[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0972_ (.CLK(clknet_4_13_0_clk),
    .D(_0024_),
    .RESET_B(_0002_),
    .Q(\top[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0973_ (.CLK(clknet_4_13_0_clk),
    .D(_0025_),
    .RESET_B(_0003_),
    .Q(\top[3] ));
 sky130_fd_sc_hd__dfrtp_2 _0974_ (.CLK(clknet_4_6_0_clk),
    .D(_0026_),
    .RESET_B(_0004_),
    .Q(\top[4] ));
 sky130_fd_sc_hd__dfrtp_1 _0975_ (.CLK(clknet_4_13_0_clk),
    .D(_0479_),
    .RESET_B(_0005_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _0976_ (.CLK(clknet_4_4_0_clk),
    .D(net31),
    .RESET_B(_0006_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _0977_ (.CLK(clknet_4_4_0_clk),
    .D(net113),
    .RESET_B(_0007_),
    .Q(net13));
 sky130_fd_sc_hd__dfrtp_1 _0978_ (.CLK(clknet_4_1_0_clk),
    .D(net37),
    .RESET_B(_0008_),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _0979_ (.CLK(clknet_4_1_0_clk),
    .D(net39),
    .RESET_B(_0009_),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _0980_ (.CLK(clknet_4_5_0_clk),
    .D(net33),
    .RESET_B(_0010_),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _0981_ (.CLK(clknet_4_3_0_clk),
    .D(net43),
    .RESET_B(_0011_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _0982_ (.CLK(clknet_4_7_0_clk),
    .D(net35),
    .RESET_B(_0012_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(clknet_4_7_0_clk),
    .D(_0034_),
    .RESET_B(_0013_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _0984_ (.CLK(clknet_4_4_0_clk),
    .D(_0035_),
    .Q(\stack[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0985_ (.CLK(clknet_4_4_0_clk),
    .D(_0036_),
    .Q(\stack[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0986_ (.CLK(clknet_4_1_0_clk),
    .D(_0037_),
    .Q(\stack[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0987_ (.CLK(clknet_4_3_0_clk),
    .D(_0038_),
    .Q(\stack[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0988_ (.CLK(clknet_4_5_0_clk),
    .D(_0039_),
    .Q(\stack[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0989_ (.CLK(clknet_4_3_0_clk),
    .D(_0040_),
    .Q(\stack[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0990_ (.CLK(clknet_4_7_0_clk),
    .D(_0041_),
    .Q(\stack[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0991_ (.CLK(clknet_4_7_0_clk),
    .D(_0042_),
    .Q(\stack[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _0992_ (.CLK(clknet_4_3_0_clk),
    .D(_0043_),
    .Q(\stack[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _0993_ (.CLK(clknet_4_1_0_clk),
    .D(_0044_),
    .Q(\stack[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _0994_ (.CLK(clknet_4_1_0_clk),
    .D(_0045_),
    .Q(\stack[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _0995_ (.CLK(clknet_4_2_0_clk),
    .D(_0046_),
    .Q(\stack[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _0996_ (.CLK(clknet_4_5_0_clk),
    .D(_0047_),
    .Q(\stack[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _0997_ (.CLK(clknet_4_2_0_clk),
    .D(_0048_),
    .Q(\stack[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _0998_ (.CLK(clknet_4_7_0_clk),
    .D(_0049_),
    .Q(\stack[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _0999_ (.CLK(clknet_4_5_0_clk),
    .D(_0050_),
    .Q(\stack[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1000_ (.CLK(clknet_4_2_0_clk),
    .D(_0051_),
    .Q(\stack[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1001_ (.CLK(clknet_4_0_0_clk),
    .D(_0052_),
    .Q(\stack[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1002_ (.CLK(clknet_4_0_0_clk),
    .D(_0053_),
    .Q(\stack[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1003_ (.CLK(clknet_4_2_0_clk),
    .D(_0054_),
    .Q(\stack[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1004_ (.CLK(clknet_4_4_0_clk),
    .D(_0055_),
    .Q(\stack[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1005_ (.CLK(clknet_4_8_0_clk),
    .D(_0056_),
    .Q(\stack[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1006_ (.CLK(clknet_4_6_0_clk),
    .D(_0057_),
    .Q(\stack[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1007_ (.CLK(clknet_4_5_0_clk),
    .D(_0058_),
    .Q(\stack[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1008_ (.CLK(clknet_4_10_0_clk),
    .D(_0059_),
    .Q(\stack[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1009_ (.CLK(clknet_4_10_0_clk),
    .D(_0060_),
    .Q(\stack[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1010_ (.CLK(clknet_4_8_0_clk),
    .D(_0061_),
    .Q(\stack[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1011_ (.CLK(clknet_4_10_0_clk),
    .D(_0062_),
    .Q(\stack[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1012_ (.CLK(clknet_4_13_0_clk),
    .D(_0063_),
    .Q(\stack[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1013_ (.CLK(clknet_4_10_0_clk),
    .D(_0064_),
    .Q(\stack[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1014_ (.CLK(clknet_4_15_0_clk),
    .D(_0065_),
    .Q(\stack[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1015_ (.CLK(clknet_4_12_0_clk),
    .D(_0066_),
    .Q(\stack[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1016_ (.CLK(clknet_4_2_0_clk),
    .D(_0067_),
    .Q(\stack[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1017_ (.CLK(clknet_4_0_0_clk),
    .D(_0068_),
    .Q(\stack[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1018_ (.CLK(clknet_4_0_0_clk),
    .D(_0069_),
    .Q(\stack[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1019_ (.CLK(clknet_4_2_0_clk),
    .D(_0070_),
    .Q(\stack[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1020_ (.CLK(clknet_4_5_0_clk),
    .D(_0071_),
    .Q(\stack[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1021_ (.CLK(clknet_4_8_0_clk),
    .D(_0072_),
    .Q(\stack[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1022_ (.CLK(clknet_4_6_0_clk),
    .D(_0073_),
    .Q(\stack[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1023_ (.CLK(clknet_4_5_0_clk),
    .D(_0074_),
    .Q(\stack[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1024_ (.CLK(clknet_4_14_0_clk),
    .D(_0075_),
    .Q(\stack[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1025_ (.CLK(clknet_4_11_0_clk),
    .D(_0076_),
    .Q(\stack[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1026_ (.CLK(clknet_4_9_0_clk),
    .D(_0077_),
    .Q(\stack[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1027_ (.CLK(clknet_4_11_0_clk),
    .D(_0078_),
    .Q(\stack[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1028_ (.CLK(clknet_4_15_0_clk),
    .D(_0079_),
    .Q(\stack[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1029_ (.CLK(clknet_4_11_0_clk),
    .D(_0080_),
    .Q(\stack[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1030_ (.CLK(clknet_4_15_0_clk),
    .D(_0081_),
    .Q(\stack[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1031_ (.CLK(clknet_4_13_0_clk),
    .D(_0082_),
    .Q(\stack[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1032_ (.CLK(clknet_4_9_0_clk),
    .D(_0083_),
    .Q(\stack[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1033_ (.CLK(clknet_4_1_0_clk),
    .D(_0084_),
    .Q(\stack[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1034_ (.CLK(clknet_4_1_0_clk),
    .D(_0085_),
    .Q(\stack[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1035_ (.CLK(clknet_4_3_0_clk),
    .D(_0086_),
    .Q(\stack[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1036_ (.CLK(clknet_4_5_0_clk),
    .D(_0087_),
    .Q(\stack[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1037_ (.CLK(clknet_4_9_0_clk),
    .D(_0088_),
    .Q(\stack[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1038_ (.CLK(clknet_4_7_0_clk),
    .D(_0089_),
    .Q(\stack[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1039_ (.CLK(clknet_4_5_0_clk),
    .D(_0090_),
    .Q(\stack[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1040_ (.CLK(clknet_4_11_0_clk),
    .D(_0091_),
    .Q(\stack[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1041_ (.CLK(clknet_4_10_0_clk),
    .D(_0092_),
    .Q(\stack[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1042_ (.CLK(clknet_4_9_0_clk),
    .D(_0093_),
    .Q(\stack[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1043_ (.CLK(clknet_4_11_0_clk),
    .D(_0094_),
    .Q(\stack[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1044_ (.CLK(clknet_4_15_0_clk),
    .D(_0095_),
    .Q(\stack[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1045_ (.CLK(clknet_4_10_0_clk),
    .D(_0096_),
    .Q(\stack[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1046_ (.CLK(clknet_4_15_0_clk),
    .D(_0097_),
    .Q(\stack[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1047_ (.CLK(clknet_4_13_0_clk),
    .D(_0098_),
    .Q(\stack[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1048_ (.CLK(clknet_4_14_0_clk),
    .D(_0099_),
    .Q(\stack[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1049_ (.CLK(clknet_4_12_0_clk),
    .D(_0100_),
    .Q(\stack[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1050_ (.CLK(clknet_4_9_0_clk),
    .D(_0101_),
    .Q(\stack[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1051_ (.CLK(clknet_4_11_0_clk),
    .D(_0102_),
    .Q(\stack[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1052_ (.CLK(clknet_4_14_0_clk),
    .D(_0103_),
    .Q(\stack[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1053_ (.CLK(clknet_4_14_0_clk),
    .D(_0104_),
    .Q(\stack[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1054_ (.CLK(clknet_4_14_0_clk),
    .D(_0105_),
    .Q(\stack[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1055_ (.CLK(clknet_4_12_0_clk),
    .D(_0106_),
    .Q(\stack[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1056_ (.CLK(clknet_4_14_0_clk),
    .D(_0107_),
    .Q(\stack[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1057_ (.CLK(clknet_4_12_0_clk),
    .D(_0108_),
    .Q(\stack[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1058_ (.CLK(clknet_4_9_0_clk),
    .D(_0109_),
    .Q(\stack[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1059_ (.CLK(clknet_4_11_0_clk),
    .D(_0110_),
    .Q(\stack[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1060_ (.CLK(clknet_4_14_0_clk),
    .D(_0111_),
    .Q(\stack[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1061_ (.CLK(clknet_4_11_0_clk),
    .D(_0112_),
    .Q(\stack[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1062_ (.CLK(clknet_4_14_0_clk),
    .D(_0113_),
    .Q(\stack[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1063_ (.CLK(clknet_4_12_0_clk),
    .D(_0114_),
    .Q(\stack[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1064_ (.CLK(clknet_4_2_0_clk),
    .D(_0115_),
    .Q(\stack[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1065_ (.CLK(clknet_4_0_0_clk),
    .D(_0116_),
    .Q(\stack[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1066_ (.CLK(clknet_4_0_0_clk),
    .D(_0117_),
    .Q(\stack[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1067_ (.CLK(clknet_4_2_0_clk),
    .D(_0118_),
    .Q(\stack[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1068_ (.CLK(clknet_4_4_0_clk),
    .D(_0119_),
    .Q(\stack[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1069_ (.CLK(clknet_4_8_0_clk),
    .D(_0120_),
    .Q(\stack[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1070_ (.CLK(clknet_4_6_0_clk),
    .D(_0121_),
    .Q(\stack[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1071_ (.CLK(clknet_4_4_0_clk),
    .D(_0122_),
    .Q(\stack[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1072_ (.CLK(clknet_4_2_0_clk),
    .D(_0123_),
    .Q(\stack[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1073_ (.CLK(clknet_4_2_0_clk),
    .D(_0124_),
    .Q(\stack[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1074_ (.CLK(clknet_4_0_0_clk),
    .D(_0125_),
    .Q(\stack[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1075_ (.CLK(clknet_4_2_0_clk),
    .D(_0126_),
    .Q(\stack[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1076_ (.CLK(clknet_4_4_0_clk),
    .D(_0127_),
    .Q(\stack[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1077_ (.CLK(clknet_4_8_0_clk),
    .D(_0128_),
    .Q(\stack[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1078_ (.CLK(clknet_4_6_0_clk),
    .D(_0129_),
    .Q(\stack[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1079_ (.CLK(clknet_4_4_0_clk),
    .D(_0130_),
    .Q(\stack[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1080_ (.CLK(clknet_4_14_0_clk),
    .D(_0131_),
    .Q(\stack[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1081_ (.CLK(clknet_4_10_0_clk),
    .D(_0132_),
    .Q(\stack[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1082_ (.CLK(clknet_4_8_0_clk),
    .D(_0133_),
    .Q(\stack[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1083_ (.CLK(clknet_4_10_0_clk),
    .D(_0134_),
    .Q(\stack[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1084_ (.CLK(clknet_4_15_0_clk),
    .D(_0135_),
    .Q(\stack[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1085_ (.CLK(clknet_4_10_0_clk),
    .D(_0136_),
    .Q(\stack[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1086_ (.CLK(clknet_4_15_0_clk),
    .D(_0137_),
    .Q(\stack[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1087_ (.CLK(clknet_4_13_0_clk),
    .D(_0138_),
    .Q(\stack[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1088_ (.CLK(clknet_4_10_0_clk),
    .D(_0139_),
    .Q(\stack[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1089_ (.CLK(clknet_4_8_0_clk),
    .D(_0140_),
    .Q(\stack[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1090_ (.CLK(clknet_4_8_0_clk),
    .D(_0141_),
    .Q(\stack[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1091_ (.CLK(clknet_4_10_0_clk),
    .D(_0142_),
    .Q(\stack[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1092_ (.CLK(clknet_4_15_0_clk),
    .D(_0143_),
    .Q(\stack[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1093_ (.CLK(clknet_4_10_0_clk),
    .D(_0144_),
    .Q(\stack[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1094_ (.CLK(clknet_4_15_0_clk),
    .D(_0145_),
    .Q(\stack[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1095_ (.CLK(clknet_4_12_0_clk),
    .D(_0146_),
    .Q(\stack[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _1096_ (.CLK(clknet_4_9_0_clk),
    .D(_0147_),
    .Q(\stack[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _1097_ (.CLK(clknet_4_1_0_clk),
    .D(_0148_),
    .Q(\stack[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _1098_ (.CLK(clknet_4_0_0_clk),
    .D(_0149_),
    .Q(\stack[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _1099_ (.CLK(clknet_4_2_0_clk),
    .D(_0150_),
    .Q(\stack[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _1100_ (.CLK(clknet_4_5_0_clk),
    .D(_0151_),
    .Q(\stack[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _1101_ (.CLK(clknet_4_9_0_clk),
    .D(_0152_),
    .Q(\stack[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _1102_ (.CLK(clknet_4_6_0_clk),
    .D(_0153_),
    .Q(\stack[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _1103_ (.CLK(clknet_4_5_0_clk),
    .D(_0154_),
    .Q(\stack[14][7] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net12),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0030_),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\stack[2][6] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\stack[15][1] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\stack[6][6] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\stack[3][4] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\stack[15][0] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\stack[9][6] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\stack[0][1] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\stack[6][2] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\stack[12][0] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\stack[6][0] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\stack[9][1] ),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\stack[10][0] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\stack[13][6] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\stack[11][3] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\stack[3][6] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\stack[14][3] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\stack[12][6] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\stack[0][4] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\stack[0][3] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\stack[15][6] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\stack[0][7] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\stack[10][6] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\stack[11][1] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\stack[3][3] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\stack[3][1] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\stack[15][7] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\stack[13][5] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\stack[3][5] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\stack[12][3] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\stack[1][5] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\stack[3][0] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\stack[12][2] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net17),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net19),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\stack[13][0] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\stack[15][4] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\stack[6][7] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\stack[1][2] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\stack[1][3] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\stack[1][4] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\stack[4][4] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\stack[6][4] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\stack[15][2] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0032_),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\stack[2][0] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\stack[1][7] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\stack[1][6] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\stack[1][1] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\stack[7][6] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\stack[9][7] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\stack[4][2] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\stack[14][6] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\stack[14][0] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0027_),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\stack[14][5] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\stack[8][1] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\stack[8][3] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\stack[8][0] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\stack[4][6] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\stack[7][2] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\stack[7][3] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\stack[13][7] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\stack[4][1] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\stack[9][3] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net16),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\stack[10][1] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\stack[13][2] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\stack[5][6] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\stack[4][5] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\stack[11][4] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\stack[14][2] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\stack[10][2] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\stack[5][5] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\stack[5][3] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\stack[11][5] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0031_),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\stack[5][1] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\stack[12][7] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\stack[5][2] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\stack[4][0] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\stack[8][7] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\stack[8][6] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\stack[8][5] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\stack[11][2] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\stack[10][5] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\stack[5][0] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net18),
    .X(net34));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\stack[7][7] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\stack[11][6] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\stack[7][0] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\stack[11][0] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\stack[7][4] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\stack[9][2] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\stack[5][7] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\stack[0][6] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\stack[2][2] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\stack[13][3] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0033_),
    .X(net35));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\stack[13][1] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\stack[14][4] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\stack[5][4] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\stack[8][2] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\stack[9][5] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\stack[10][4] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\stack[2][4] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\stack[3][7] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\stack[2][7] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\stack[14][1] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net14),
    .X(net36));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\stack[12][1] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\stack[9][0] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\stack[6][5] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\stack[7][1] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\stack[0][2] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\stack[2][3] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\stack[10][7] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\stack[0][5] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\stack[2][5] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\stack[8][4] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0029_),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\stack[1][0] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\stack[6][3] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\stack[15][5] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net13),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0028_),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\stack[11][7] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\stack[4][3] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\stack[12][4] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\stack[4][7] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\stack[15][3] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net15),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\stack[2][1] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\stack[3][2] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\stack[13][4] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\stack[0][0] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\stack[6][1] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\stack[7][5] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\stack[9][4] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\stack[10][3] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\stack[12][5] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\stack[14][7] ),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(push),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(data_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(data_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(data_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(data_in[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(data_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(data_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(data_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(pop),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap24 (.A(_0193_),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 max_cap25 (.A(_0191_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 max_cap26 (.A(_0191_),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 max_cap28 (.A(net173),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 max_cap29 (.A(_0158_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_4 output13 (.A(net13),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output14 (.A(net14),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_4 output15 (.A(net15),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_4 output17 (.A(net17),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_4 output18 (.A(net18),
    .X(data_out[6]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_4 output20 (.A(net20),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_4 output21 (.A(net21),
    .X(error));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(full));
 sky130_fd_sc_hd__buf_1 wire1 (.A(_0183_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 wire23 (.A(_0193_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 wire27 (.A(net173),
    .X(net27));
endmodule

