magic
tech sky130A
magscale 1 2
timestamp 1755431346
<< checkpaint >>
rect -1260 8876 33712 35856
rect -2590 372 33712 8876
rect -1260 -1260 33712 372
<< viali >>
rect 17877 31977 17911 32011
rect 24593 31977 24627 32011
rect 7573 31909 7607 31943
rect 1501 31773 1535 31807
rect 1685 31773 1719 31807
rect 7297 31773 7331 31807
rect 12357 31773 12391 31807
rect 18153 31773 18187 31807
rect 18889 31773 18923 31807
rect 24501 31773 24535 31807
rect 29745 31773 29779 31807
rect 12541 31637 12575 31671
rect 18337 31637 18371 31671
rect 29929 31637 29963 31671
rect 11529 31433 11563 31467
rect 17969 31433 18003 31467
rect 18061 31365 18095 31399
rect 11161 31297 11195 31331
rect 11897 31297 11931 31331
rect 12357 31297 12391 31331
rect 18797 31297 18831 31331
rect 19257 31297 19291 31331
rect 20729 31297 20763 31331
rect 21373 31297 21407 31331
rect 23857 31297 23891 31331
rect 7665 31229 7699 31263
rect 11989 31229 12023 31263
rect 12173 31229 12207 31263
rect 12909 31229 12943 31263
rect 18153 31229 18187 31263
rect 18889 31229 18923 31263
rect 18981 31229 19015 31263
rect 19809 31229 19843 31263
rect 22385 31229 22419 31263
rect 23305 31229 23339 31263
rect 24685 31229 24719 31263
rect 18429 31161 18463 31195
rect 7021 31093 7055 31127
rect 10977 31093 11011 31127
rect 17601 31093 17635 31127
rect 20545 31093 20579 31127
rect 21557 31093 21591 31127
rect 21833 31093 21867 31127
rect 22753 31093 22787 31127
rect 24041 31093 24075 31127
rect 24133 31093 24167 31127
rect 12081 30889 12115 30923
rect 18705 30889 18739 30923
rect 23121 30889 23155 30923
rect 24225 30889 24259 30923
rect 24409 30889 24443 30923
rect 9597 30753 9631 30787
rect 10701 30753 10735 30787
rect 13553 30753 13587 30787
rect 23673 30753 23707 30787
rect 5457 30685 5491 30719
rect 5733 30685 5767 30719
rect 7389 30685 7423 30719
rect 10333 30685 10367 30719
rect 10968 30685 11002 30719
rect 13737 30685 13771 30719
rect 14105 30685 14139 30719
rect 16129 30685 16163 30719
rect 16773 30685 16807 30719
rect 17049 30685 17083 30719
rect 17325 30685 17359 30719
rect 20269 30685 20303 30719
rect 21741 30685 21775 30719
rect 21997 30685 22031 30719
rect 23857 30685 23891 30719
rect 25789 30685 25823 30719
rect 5978 30617 6012 30651
rect 7656 30617 7690 30651
rect 9321 30617 9355 30651
rect 9781 30617 9815 30651
rect 13286 30617 13320 30651
rect 14350 30617 14384 30651
rect 17570 30617 17604 30651
rect 20536 30617 20570 30651
rect 25522 30617 25556 30651
rect 5641 30549 5675 30583
rect 7113 30549 7147 30583
rect 8769 30549 8803 30583
rect 8953 30549 8987 30583
rect 9413 30549 9447 30583
rect 12173 30549 12207 30583
rect 13921 30549 13955 30583
rect 15485 30549 15519 30583
rect 15577 30549 15611 30583
rect 16957 30549 16991 30583
rect 17233 30549 17267 30583
rect 21649 30549 21683 30583
rect 23765 30549 23799 30583
rect 6377 30345 6411 30379
rect 8125 30345 8159 30379
rect 14013 30345 14047 30379
rect 20637 30345 20671 30379
rect 21005 30345 21039 30379
rect 22201 30345 22235 30379
rect 6745 30277 6779 30311
rect 11897 30277 11931 30311
rect 11989 30277 12023 30311
rect 14381 30277 14415 30311
rect 1409 30209 1443 30243
rect 8309 30209 8343 30243
rect 10977 30209 11011 30243
rect 12357 30209 12391 30243
rect 12909 30209 12943 30243
rect 17233 30209 17267 30243
rect 17489 30209 17523 30243
rect 21097 30209 21131 30243
rect 22293 30209 22327 30243
rect 23029 30209 23063 30243
rect 23305 30209 23339 30243
rect 23561 30209 23595 30243
rect 6837 30141 6871 30175
rect 6929 30141 6963 30175
rect 12081 30141 12115 30175
rect 14473 30141 14507 30175
rect 14565 30141 14599 30175
rect 21281 30141 21315 30175
rect 22477 30141 22511 30175
rect 25329 30141 25363 30175
rect 1593 30073 1627 30107
rect 11529 30073 11563 30107
rect 18613 30073 18647 30107
rect 23213 30073 23247 30107
rect 11161 30005 11195 30039
rect 21833 30005 21867 30039
rect 24685 30005 24719 30039
rect 24777 30005 24811 30039
rect 23489 29801 23523 29835
rect 19993 29733 20027 29767
rect 24133 29665 24167 29699
rect 8493 29597 8527 29631
rect 9965 29597 9999 29631
rect 10149 29597 10183 29631
rect 10425 29597 10459 29631
rect 10517 29597 10551 29631
rect 12357 29597 12391 29631
rect 14657 29597 14691 29631
rect 16681 29597 16715 29631
rect 19441 29597 19475 29631
rect 19717 29597 19751 29631
rect 19809 29597 19843 29631
rect 21005 29597 21039 29631
rect 22845 29597 22879 29631
rect 23029 29597 23063 29631
rect 23121 29597 23155 29631
rect 23213 29597 23247 29631
rect 23857 29597 23891 29631
rect 25973 29597 26007 29631
rect 10333 29529 10367 29563
rect 14924 29529 14958 29563
rect 19625 29529 19659 29563
rect 25728 29529 25762 29563
rect 8309 29461 8343 29495
rect 9413 29461 9447 29495
rect 10701 29461 10735 29495
rect 11713 29461 11747 29495
rect 16037 29461 16071 29495
rect 16129 29461 16163 29495
rect 20821 29461 20855 29495
rect 23397 29461 23431 29495
rect 23949 29461 23983 29495
rect 24593 29461 24627 29495
rect 9321 29257 9355 29291
rect 11897 29257 11931 29291
rect 14473 29257 14507 29291
rect 14841 29257 14875 29291
rect 15025 29257 15059 29291
rect 15393 29257 15427 29291
rect 17969 29257 18003 29291
rect 20085 29257 20119 29291
rect 26249 29257 26283 29291
rect 8208 29189 8242 29223
rect 12633 29189 12667 29223
rect 15485 29189 15519 29223
rect 18429 29189 18463 29223
rect 19717 29189 19751 29223
rect 20536 29189 20570 29223
rect 24317 29189 24351 29223
rect 6561 29121 6595 29155
rect 7941 29121 7975 29155
rect 10232 29121 10266 29155
rect 12541 29121 12575 29155
rect 12725 29121 12759 29155
rect 12909 29121 12943 29155
rect 13093 29121 13127 29155
rect 13349 29121 13383 29155
rect 14657 29121 14691 29155
rect 17877 29121 17911 29155
rect 18337 29121 18371 29155
rect 18797 29121 18831 29155
rect 19533 29121 19567 29155
rect 19809 29121 19843 29155
rect 19901 29121 19935 29155
rect 24225 29121 24259 29155
rect 24409 29121 24443 29155
rect 24593 29121 24627 29155
rect 25053 29121 25087 29155
rect 25513 29121 25547 29155
rect 26065 29121 26099 29155
rect 26433 29121 26467 29155
rect 6101 29053 6135 29087
rect 9965 29053 9999 29087
rect 11989 29053 12023 29087
rect 12173 29053 12207 29087
rect 15669 29053 15703 29087
rect 18613 29053 18647 29087
rect 19349 29053 19383 29087
rect 20269 29053 20303 29087
rect 22477 29053 22511 29087
rect 24777 29053 24811 29087
rect 24961 29053 24995 29087
rect 11345 28985 11379 29019
rect 21649 28985 21683 29019
rect 25421 28985 25455 29019
rect 5549 28917 5583 28951
rect 6377 28917 6411 28951
rect 11529 28917 11563 28951
rect 12357 28917 12391 28951
rect 17693 28917 17727 28951
rect 21833 28917 21867 28951
rect 24041 28917 24075 28951
rect 7021 28713 7055 28747
rect 8953 28713 8987 28747
rect 10517 28713 10551 28747
rect 13001 28713 13035 28747
rect 15485 28713 15519 28747
rect 15577 28713 15611 28747
rect 18797 28713 18831 28747
rect 20821 28713 20855 28747
rect 6929 28645 6963 28679
rect 12633 28645 12667 28679
rect 7573 28577 7607 28611
rect 8401 28577 8435 28611
rect 9597 28577 9631 28611
rect 13553 28577 13587 28611
rect 13737 28577 13771 28611
rect 14657 28577 14691 28611
rect 19809 28577 19843 28611
rect 20729 28577 20763 28611
rect 21373 28577 21407 28611
rect 5549 28509 5583 28543
rect 9321 28509 9355 28543
rect 10701 28509 10735 28543
rect 12081 28509 12115 28543
rect 12357 28509 12391 28543
rect 12449 28509 12483 28543
rect 12817 28509 12851 28543
rect 14933 28509 14967 28543
rect 15117 28509 15151 28543
rect 15209 28509 15243 28543
rect 15301 28509 15335 28543
rect 15761 28509 15795 28543
rect 15853 28509 15887 28543
rect 17417 28509 17451 28543
rect 21189 28509 21223 28543
rect 5816 28441 5850 28475
rect 12265 28441 12299 28475
rect 13461 28441 13495 28475
rect 14105 28441 14139 28475
rect 15577 28441 15611 28475
rect 17662 28441 17696 28475
rect 19625 28441 19659 28475
rect 20085 28441 20119 28475
rect 7389 28373 7423 28407
rect 7481 28373 7515 28407
rect 7849 28373 7883 28407
rect 9413 28373 9447 28407
rect 13093 28373 13127 28407
rect 16037 28373 16071 28407
rect 19257 28373 19291 28407
rect 19717 28373 19751 28407
rect 21281 28373 21315 28407
rect 5733 28169 5767 28203
rect 5825 28169 5859 28203
rect 9137 28169 9171 28203
rect 17417 28169 17451 28203
rect 22385 28169 22419 28203
rect 8861 28101 8895 28135
rect 12817 28101 12851 28135
rect 23581 28101 23615 28135
rect 3893 28033 3927 28067
rect 4160 28033 4194 28067
rect 6377 28033 6411 28067
rect 6633 28033 6667 28067
rect 8585 28033 8619 28067
rect 8769 28033 8803 28067
rect 8953 28033 8987 28067
rect 10701 28033 10735 28067
rect 10977 28033 11011 28067
rect 12633 28033 12667 28067
rect 12909 28033 12943 28067
rect 17233 28033 17267 28067
rect 17776 28033 17810 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22109 28033 22143 28067
rect 22201 28033 22235 28067
rect 22937 28033 22971 28067
rect 23213 28033 23247 28067
rect 23857 28033 23891 28067
rect 6009 27965 6043 27999
rect 8401 27965 8435 27999
rect 10885 27965 10919 27999
rect 12449 27965 12483 27999
rect 17509 27965 17543 27999
rect 23029 27965 23063 27999
rect 23765 27965 23799 27999
rect 5273 27897 5307 27931
rect 7757 27897 7791 27931
rect 18889 27897 18923 27931
rect 5365 27829 5399 27863
rect 7849 27829 7883 27863
rect 10977 27829 11011 27863
rect 11161 27829 11195 27863
rect 22937 27829 22971 27863
rect 23397 27829 23431 27863
rect 23581 27829 23615 27863
rect 24041 27829 24075 27863
rect 4261 27625 4295 27659
rect 6101 27625 6135 27659
rect 13645 27625 13679 27659
rect 16405 27625 16439 27659
rect 22017 27625 22051 27659
rect 23397 27625 23431 27659
rect 6193 27557 6227 27591
rect 7573 27557 7607 27591
rect 6837 27489 6871 27523
rect 14657 27489 14691 27523
rect 21005 27489 21039 27523
rect 21373 27489 21407 27523
rect 22753 27489 22787 27523
rect 24869 27489 24903 27523
rect 4445 27421 4479 27455
rect 5917 27421 5951 27455
rect 6653 27421 6687 27455
rect 7021 27421 7055 27455
rect 7205 27421 7239 27455
rect 7389 27421 7423 27455
rect 11989 27421 12023 27455
rect 12265 27421 12299 27455
rect 15761 27421 15795 27455
rect 16589 27421 16623 27455
rect 16865 27421 16899 27455
rect 17141 27421 17175 27455
rect 20821 27421 20855 27455
rect 21557 27421 21591 27455
rect 22845 27421 22879 27455
rect 23213 27421 23247 27455
rect 25053 27421 25087 27455
rect 26157 27421 26191 27455
rect 7297 27353 7331 27387
rect 12510 27353 12544 27387
rect 20913 27353 20947 27387
rect 22109 27353 22143 27387
rect 23029 27353 23063 27387
rect 23121 27353 23155 27387
rect 25145 27353 25179 27387
rect 25605 27353 25639 27387
rect 26709 27353 26743 27387
rect 6561 27285 6595 27319
rect 12173 27285 12207 27319
rect 14105 27285 14139 27319
rect 16313 27285 16347 27319
rect 16773 27285 16807 27319
rect 16957 27285 16991 27319
rect 20453 27285 20487 27319
rect 21649 27285 21683 27319
rect 25513 27285 25547 27319
rect 26617 27285 26651 27319
rect 12725 27081 12759 27115
rect 13093 27081 13127 27115
rect 15117 27081 15151 27115
rect 19993 27081 20027 27115
rect 21833 27081 21867 27115
rect 23581 27081 23615 27115
rect 24133 27081 24167 27115
rect 24501 27081 24535 27115
rect 24777 27081 24811 27115
rect 26249 27081 26283 27115
rect 13185 27013 13219 27047
rect 16252 27013 16286 27047
rect 20330 27013 20364 27047
rect 23949 27013 23983 27047
rect 25912 27013 25946 27047
rect 19809 26945 19843 26979
rect 22753 26945 22787 26979
rect 23765 26945 23799 26979
rect 24041 26945 24075 26979
rect 24317 26945 24351 26979
rect 24593 26945 24627 26979
rect 26157 26945 26191 26979
rect 26433 26945 26467 26979
rect 10701 26877 10735 26911
rect 13369 26877 13403 26911
rect 16497 26877 16531 26911
rect 20085 26877 20119 26911
rect 22477 26877 22511 26911
rect 21465 26809 21499 26843
rect 10057 26741 10091 26775
rect 22569 26741 22603 26775
rect 16497 26537 16531 26571
rect 18981 26537 19015 26571
rect 21833 26537 21867 26571
rect 10333 26469 10367 26503
rect 25789 26469 25823 26503
rect 13737 26401 13771 26435
rect 15945 26401 15979 26435
rect 17049 26401 17083 26435
rect 24409 26401 24443 26435
rect 8585 26333 8619 26367
rect 8953 26333 8987 26367
rect 11069 26333 11103 26367
rect 11161 26333 11195 26367
rect 11437 26333 11471 26367
rect 11529 26333 11563 26367
rect 13553 26333 13587 26367
rect 14657 26333 14691 26367
rect 16129 26333 16163 26367
rect 18705 26333 18739 26367
rect 20453 26333 20487 26367
rect 24041 26333 24075 26367
rect 9198 26265 9232 26299
rect 11345 26265 11379 26299
rect 13461 26265 13495 26299
rect 14105 26265 14139 26299
rect 16037 26265 16071 26299
rect 17877 26265 17911 26299
rect 20720 26265 20754 26299
rect 24654 26265 24688 26299
rect 8769 26197 8803 26231
rect 10425 26197 10459 26231
rect 11713 26197 11747 26231
rect 13093 26197 13127 26231
rect 24225 26197 24259 26231
rect 9321 25993 9355 26027
rect 9689 25993 9723 26027
rect 10517 25993 10551 26027
rect 12817 25993 12851 26027
rect 14289 25993 14323 26027
rect 24225 25993 24259 26027
rect 10609 25925 10643 25959
rect 13176 25925 13210 25959
rect 19993 25925 20027 25959
rect 7849 25857 7883 25891
rect 8116 25857 8150 25891
rect 9781 25857 9815 25891
rect 12633 25857 12667 25891
rect 19165 25857 19199 25891
rect 24593 25857 24627 25891
rect 25053 25857 25087 25891
rect 25697 25857 25731 25891
rect 5549 25789 5583 25823
rect 9965 25789 9999 25823
rect 10701 25789 10735 25823
rect 12909 25789 12943 25823
rect 24685 25789 24719 25823
rect 24777 25789 24811 25823
rect 9229 25721 9263 25755
rect 4905 25653 4939 25687
rect 10149 25653 10183 25687
rect 8217 25449 8251 25483
rect 30849 25449 30883 25483
rect 6469 25381 6503 25415
rect 10977 25381 11011 25415
rect 4905 25313 4939 25347
rect 7205 25313 7239 25347
rect 7941 25313 7975 25347
rect 9597 25313 9631 25347
rect 11621 25313 11655 25347
rect 18061 25313 18095 25347
rect 18889 25313 18923 25347
rect 4169 25245 4203 25279
rect 4629 25245 4663 25279
rect 5089 25245 5123 25279
rect 8401 25245 8435 25279
rect 9321 25245 9355 25279
rect 12081 25245 12115 25279
rect 14749 25245 14783 25279
rect 17969 25245 18003 25279
rect 19809 25245 19843 25279
rect 30665 25245 30699 25279
rect 5356 25177 5390 25211
rect 9842 25177 9876 25211
rect 12348 25177 12382 25211
rect 17877 25177 17911 25211
rect 18705 25177 18739 25211
rect 19257 25177 19291 25211
rect 3985 25109 4019 25143
rect 4261 25109 4295 25143
rect 4721 25109 4755 25143
rect 6561 25109 6595 25143
rect 6929 25109 6963 25143
rect 7021 25109 7055 25143
rect 7389 25109 7423 25143
rect 9505 25109 9539 25143
rect 11069 25109 11103 25143
rect 13461 25109 13495 25143
rect 14105 25109 14139 25143
rect 17509 25109 17543 25143
rect 18337 25109 18371 25143
rect 18797 25109 18831 25143
rect 5457 24905 5491 24939
rect 9597 24905 9631 24939
rect 9965 24905 9999 24939
rect 12265 24905 12299 24939
rect 12909 24905 12943 24939
rect 18981 24905 19015 24939
rect 6653 24837 6687 24871
rect 8125 24837 8159 24871
rect 11253 24837 11287 24871
rect 20729 24837 20763 24871
rect 21833 24837 21867 24871
rect 3709 24769 3743 24803
rect 3976 24769 4010 24803
rect 5641 24769 5675 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6745 24769 6779 24803
rect 8953 24769 8987 24803
rect 10425 24769 10459 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 11805 24769 11839 24803
rect 11897 24769 11931 24803
rect 12449 24769 12483 24803
rect 13001 24769 13035 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 13829 24769 13863 24803
rect 17417 24769 17451 24803
rect 17765 24769 17799 24803
rect 19717 24769 19751 24803
rect 19901 24769 19935 24803
rect 19993 24769 20027 24803
rect 20085 24769 20119 24803
rect 20821 24769 20855 24803
rect 21373 24769 21407 24803
rect 10057 24701 10091 24735
rect 10149 24701 10183 24735
rect 13185 24701 13219 24735
rect 14933 24701 14967 24735
rect 17509 24701 17543 24735
rect 19533 24701 19567 24735
rect 20913 24701 20947 24735
rect 22385 24701 22419 24735
rect 24409 24701 24443 24735
rect 25237 24701 25271 24735
rect 5089 24633 5123 24667
rect 12541 24633 12575 24667
rect 20361 24633 20395 24667
rect 6929 24565 6963 24599
rect 12081 24565 12115 24599
rect 13369 24565 13403 24599
rect 14381 24565 14415 24599
rect 17233 24565 17267 24599
rect 18889 24565 18923 24599
rect 20269 24565 20303 24599
rect 21189 24565 21223 24599
rect 23857 24565 23891 24599
rect 24593 24565 24627 24599
rect 11989 24361 12023 24395
rect 14289 24361 14323 24395
rect 18429 24361 18463 24395
rect 21281 24361 21315 24395
rect 21373 24361 21407 24395
rect 24041 24361 24075 24395
rect 11897 24225 11931 24259
rect 15669 24225 15703 24259
rect 21925 24225 21959 24259
rect 24961 24225 24995 24259
rect 25329 24225 25363 24259
rect 8585 24157 8619 24191
rect 10333 24157 10367 24191
rect 11713 24157 11747 24191
rect 11989 24157 12023 24191
rect 16313 24157 16347 24191
rect 17049 24157 17083 24191
rect 17316 24157 17350 24191
rect 19625 24157 19659 24191
rect 19901 24157 19935 24191
rect 21741 24157 21775 24191
rect 22661 24157 22695 24191
rect 24777 24157 24811 24191
rect 1501 24089 1535 24123
rect 1869 24089 1903 24123
rect 15402 24089 15436 24123
rect 20157 24089 20191 24123
rect 22928 24089 22962 24123
rect 24869 24089 24903 24123
rect 25513 24089 25547 24123
rect 8401 24021 8435 24055
rect 9689 24021 9723 24055
rect 11529 24021 11563 24055
rect 15761 24021 15795 24055
rect 19809 24021 19843 24055
rect 21833 24021 21867 24055
rect 24409 24021 24443 24055
rect 25605 24021 25639 24055
rect 25973 24021 26007 24055
rect 9505 23817 9539 23851
rect 9873 23817 9907 23851
rect 13829 23817 13863 23851
rect 13921 23817 13955 23851
rect 14289 23817 14323 23851
rect 14749 23817 14783 23851
rect 17601 23817 17635 23851
rect 21833 23817 21867 23851
rect 23489 23817 23523 23851
rect 24225 23817 24259 23851
rect 25789 23817 25823 23851
rect 8300 23749 8334 23783
rect 17877 23749 17911 23783
rect 20352 23749 20386 23783
rect 22569 23749 22603 23783
rect 24562 23749 24596 23783
rect 4997 23681 5031 23715
rect 5457 23681 5491 23715
rect 8033 23681 8067 23715
rect 9965 23681 9999 23715
rect 12817 23681 12851 23715
rect 13001 23681 13035 23715
rect 13093 23681 13127 23715
rect 13645 23681 13679 23715
rect 15873 23681 15907 23715
rect 16129 23681 16163 23715
rect 16405 23681 16439 23715
rect 17417 23681 17451 23715
rect 18705 23681 18739 23715
rect 20085 23681 20119 23715
rect 22845 23681 22879 23715
rect 23581 23681 23615 23715
rect 24041 23681 24075 23715
rect 26709 23681 26743 23715
rect 5089 23613 5123 23647
rect 5273 23613 5307 23647
rect 6009 23613 6043 23647
rect 10057 23613 10091 23647
rect 14381 23613 14415 23647
rect 14565 23613 14599 23647
rect 22385 23613 22419 23647
rect 22753 23613 22787 23647
rect 23673 23613 23707 23647
rect 24317 23613 24351 23647
rect 26341 23613 26375 23647
rect 9413 23545 9447 23579
rect 16221 23545 16255 23579
rect 21465 23545 21499 23579
rect 4629 23477 4663 23511
rect 12633 23477 12667 23511
rect 22569 23477 22603 23511
rect 23029 23477 23063 23511
rect 23121 23477 23155 23511
rect 25697 23477 25731 23511
rect 26525 23477 26559 23511
rect 11805 23273 11839 23307
rect 13921 23273 13955 23307
rect 15761 23273 15795 23307
rect 22385 23273 22419 23307
rect 22937 23273 22971 23307
rect 23673 23273 23707 23307
rect 24501 23273 24535 23307
rect 8769 23205 8803 23239
rect 4813 23137 4847 23171
rect 6837 23137 6871 23171
rect 9413 23137 9447 23171
rect 9597 23137 9631 23171
rect 10333 23137 10367 23171
rect 11805 23137 11839 23171
rect 12541 23137 12575 23171
rect 14657 23137 14691 23171
rect 15209 23137 15243 23171
rect 21189 23137 21223 23171
rect 4445 23069 4479 23103
rect 6653 23069 6687 23103
rect 7389 23069 7423 23103
rect 10517 23069 10551 23103
rect 10701 23069 10735 23103
rect 10793 23069 10827 23103
rect 10885 23069 10919 23103
rect 11897 23069 11931 23103
rect 12265 23069 12299 23103
rect 15301 23069 15335 23103
rect 15393 23069 15427 23103
rect 21833 23069 21867 23103
rect 22109 23069 22143 23103
rect 22201 23069 22235 23103
rect 23121 23069 23155 23103
rect 23857 23069 23891 23103
rect 23949 23069 23983 23103
rect 24225 23069 24259 23103
rect 25881 23069 25915 23103
rect 5080 23001 5114 23035
rect 7656 23001 7690 23035
rect 9321 23001 9355 23035
rect 9781 23001 9815 23035
rect 11621 23001 11655 23035
rect 12786 23001 12820 23035
rect 20453 23001 20487 23035
rect 22017 23001 22051 23035
rect 24041 23001 24075 23035
rect 25636 23001 25670 23035
rect 4261 22933 4295 22967
rect 6193 22933 6227 22967
rect 6285 22933 6319 22967
rect 6745 22933 6779 22967
rect 8953 22933 8987 22967
rect 11069 22933 11103 22967
rect 12081 22933 12115 22967
rect 12449 22933 12483 22967
rect 14105 22933 14139 22967
rect 5365 22729 5399 22763
rect 6469 22729 6503 22763
rect 7849 22729 7883 22763
rect 13001 22729 13035 22763
rect 13369 22729 13403 22763
rect 14381 22729 14415 22763
rect 23765 22729 23799 22763
rect 24133 22729 24167 22763
rect 4160 22661 4194 22695
rect 7389 22661 7423 22695
rect 14657 22661 14691 22695
rect 14749 22661 14783 22695
rect 5549 22593 5583 22627
rect 7205 22593 7239 22627
rect 7481 22593 7515 22627
rect 7573 22593 7607 22627
rect 8033 22593 8067 22627
rect 13461 22593 13495 22627
rect 14565 22593 14599 22627
rect 14933 22593 14967 22627
rect 23949 22593 23983 22627
rect 24225 22593 24259 22627
rect 3893 22525 3927 22559
rect 7021 22525 7055 22559
rect 13645 22525 13679 22559
rect 5273 22457 5307 22491
rect 7757 22457 7791 22491
rect 14105 22117 14139 22151
rect 24409 22117 24443 22151
rect 8309 22049 8343 22083
rect 8493 22049 8527 22083
rect 17417 22049 17451 22083
rect 17969 22049 18003 22083
rect 19257 22049 19291 22083
rect 9321 21981 9355 22015
rect 11069 21981 11103 22015
rect 14657 21981 14691 22015
rect 15577 21981 15611 22015
rect 16773 21981 16807 22015
rect 16957 21981 16991 22015
rect 17325 21981 17359 22015
rect 23765 21981 23799 22015
rect 15393 21913 15427 21947
rect 16037 21913 16071 21947
rect 16221 21913 16255 21947
rect 16313 21913 16347 21947
rect 16497 21913 16531 21947
rect 16681 21913 16715 21947
rect 19533 21913 19567 21947
rect 24593 21913 24627 21947
rect 7849 21845 7883 21879
rect 8217 21845 8251 21879
rect 9505 21845 9539 21879
rect 10425 21845 10459 21879
rect 15853 21845 15887 21879
rect 21005 21845 21039 21879
rect 23949 21845 23983 21879
rect 8861 21641 8895 21675
rect 13093 21641 13127 21675
rect 13553 21641 13587 21675
rect 6561 21573 6595 21607
rect 8769 21573 8803 21607
rect 15301 21573 15335 21607
rect 16865 21573 16899 21607
rect 17049 21573 17083 21607
rect 21833 21573 21867 21607
rect 6377 21505 6411 21539
rect 6653 21505 6687 21539
rect 6745 21505 6779 21539
rect 9597 21505 9631 21539
rect 9853 21505 9887 21539
rect 11980 21505 12014 21539
rect 15945 21505 15979 21539
rect 16313 21505 16347 21539
rect 17325 21505 17359 21539
rect 17693 21505 17727 21539
rect 22201 21505 22235 21539
rect 23397 21505 23431 21539
rect 23765 21505 23799 21539
rect 24225 21505 24259 21539
rect 6009 21437 6043 21471
rect 7941 21437 7975 21471
rect 9505 21437 9539 21471
rect 11713 21437 11747 21471
rect 13645 21437 13679 21471
rect 13829 21437 13863 21471
rect 15853 21437 15887 21471
rect 16497 21437 16531 21471
rect 17463 21437 17497 21471
rect 17785 21437 17819 21471
rect 18061 21437 18095 21471
rect 23673 21437 23707 21471
rect 23882 21437 23916 21471
rect 16681 21369 16715 21403
rect 5457 21301 5491 21335
rect 6929 21301 6963 21335
rect 10977 21301 11011 21335
rect 13185 21301 13219 21335
rect 24041 21301 24075 21335
rect 24317 21301 24351 21335
rect 5181 21097 5215 21131
rect 8401 21097 8435 21131
rect 9413 21097 9447 21131
rect 12541 21097 12575 21131
rect 19533 21097 19567 21131
rect 20177 21097 20211 21131
rect 22385 21097 22419 21131
rect 23673 21097 23707 21131
rect 24501 21097 24535 21131
rect 5917 20961 5951 20995
rect 6377 20961 6411 20995
rect 9873 20961 9907 20995
rect 10057 20961 10091 20995
rect 15393 20961 15427 20995
rect 16129 20961 16163 20995
rect 16773 20961 16807 20995
rect 17417 20961 17451 20995
rect 17877 20961 17911 20995
rect 20729 20961 20763 20995
rect 22226 20961 22260 20995
rect 3801 20893 3835 20927
rect 5641 20893 5675 20927
rect 7021 20893 7055 20927
rect 8769 20893 8803 20927
rect 9781 20893 9815 20927
rect 10241 20893 10275 20927
rect 11621 20893 11655 20927
rect 11897 20893 11931 20927
rect 11989 20893 12023 20927
rect 12449 20893 12483 20927
rect 12725 20893 12759 20927
rect 14657 20893 14691 20927
rect 16037 20893 16071 20927
rect 16405 20893 16439 20927
rect 16589 20893 16623 20927
rect 17325 20893 17359 20927
rect 17693 20893 17727 20927
rect 18429 20893 18463 20927
rect 20085 20893 20119 20927
rect 20637 20893 20671 20927
rect 21097 20893 21131 20927
rect 21649 20893 21683 20927
rect 21741 20893 21775 20927
rect 22017 20893 22051 20927
rect 23029 20893 23063 20927
rect 23857 20893 23891 20927
rect 23949 20893 23983 20927
rect 24041 20893 24075 20927
rect 24133 20893 24167 20927
rect 4068 20825 4102 20859
rect 7288 20825 7322 20859
rect 10977 20825 11011 20859
rect 11805 20825 11839 20859
rect 17969 20825 18003 20859
rect 18153 20825 18187 20859
rect 18337 20825 18371 20859
rect 19441 20825 19475 20859
rect 21189 20825 21223 20859
rect 24593 20825 24627 20859
rect 5273 20757 5307 20791
rect 5733 20757 5767 20791
rect 6929 20757 6963 20791
rect 8585 20757 8619 20791
rect 12173 20757 12207 20791
rect 12265 20757 12299 20791
rect 14105 20757 14139 20791
rect 18613 20757 18647 20791
rect 22109 20757 22143 20791
rect 22937 20757 22971 20791
rect 4169 20553 4203 20587
rect 6193 20553 6227 20587
rect 6837 20553 6871 20587
rect 7481 20553 7515 20587
rect 9597 20553 9631 20587
rect 9689 20553 9723 20587
rect 13369 20553 13403 20587
rect 13737 20553 13771 20587
rect 15945 20553 15979 20587
rect 18337 20553 18371 20587
rect 24961 20553 24995 20587
rect 14381 20485 14415 20519
rect 16313 20485 16347 20519
rect 17049 20485 17083 20519
rect 18245 20485 18279 20519
rect 18500 20485 18534 20519
rect 18705 20485 18739 20519
rect 20729 20485 20763 20519
rect 21189 20485 21223 20519
rect 23765 20485 23799 20519
rect 25145 20485 25179 20519
rect 4353 20417 4387 20451
rect 5080 20417 5114 20451
rect 6745 20417 6779 20451
rect 7665 20417 7699 20451
rect 8217 20417 8251 20451
rect 8484 20417 8518 20451
rect 10057 20417 10091 20451
rect 10517 20417 10551 20451
rect 11069 20417 11103 20451
rect 11897 20417 11931 20451
rect 12164 20417 12198 20451
rect 15485 20417 15519 20451
rect 15669 20417 15703 20451
rect 16129 20417 16163 20451
rect 17785 20417 17819 20451
rect 18061 20417 18095 20451
rect 20637 20417 20671 20451
rect 21097 20417 21131 20451
rect 22017 20417 22051 20451
rect 22385 20417 22419 20451
rect 22569 20417 22603 20451
rect 23029 20417 23063 20451
rect 23673 20417 23707 20451
rect 24593 20417 24627 20451
rect 24685 20417 24719 20451
rect 4813 20349 4847 20383
rect 6929 20349 6963 20383
rect 10149 20349 10183 20383
rect 10333 20349 10367 20383
rect 13829 20349 13863 20383
rect 13921 20349 13955 20383
rect 14197 20349 14231 20383
rect 21649 20349 21683 20383
rect 22293 20349 22327 20383
rect 23213 20349 23247 20383
rect 23305 20349 23339 20383
rect 24225 20349 24259 20383
rect 24317 20349 24351 20383
rect 24802 20349 24836 20383
rect 13277 20281 13311 20315
rect 6377 20213 6411 20247
rect 15853 20213 15887 20247
rect 17877 20213 17911 20247
rect 18521 20213 18555 20247
rect 25237 20213 25271 20247
rect 5549 20009 5583 20043
rect 11437 20009 11471 20043
rect 18889 20009 18923 20043
rect 19257 20009 19291 20043
rect 22293 20009 22327 20043
rect 11069 19941 11103 19975
rect 19073 19941 19107 19975
rect 11345 19873 11379 19907
rect 12357 19873 12391 19907
rect 21624 19873 21658 19907
rect 23397 19873 23431 19907
rect 5733 19805 5767 19839
rect 10517 19805 10551 19839
rect 10701 19805 10735 19839
rect 10793 19805 10827 19839
rect 10885 19805 10919 19839
rect 11437 19805 11471 19839
rect 12541 19805 12575 19839
rect 12817 19805 12851 19839
rect 15945 19805 15979 19839
rect 16313 19805 16347 19839
rect 16681 19805 16715 19839
rect 19441 19805 19475 19839
rect 19717 19805 19751 19839
rect 20821 19805 20855 19839
rect 21373 19805 21407 19839
rect 22109 19805 22143 19839
rect 22385 19805 22419 19839
rect 22753 19805 22787 19839
rect 23121 19805 23155 19839
rect 23581 19805 23615 19839
rect 23857 19805 23891 19839
rect 23949 19805 23983 19839
rect 24409 19805 24443 19839
rect 26709 19805 26743 19839
rect 11161 19737 11195 19771
rect 12725 19737 12759 19771
rect 18705 19737 18739 19771
rect 20361 19737 20395 19771
rect 20453 19737 20487 19771
rect 20913 19737 20947 19771
rect 11621 19669 11655 19703
rect 18915 19669 18949 19703
rect 19625 19669 19659 19703
rect 21465 19669 21499 19703
rect 21741 19669 21775 19703
rect 21833 19669 21867 19703
rect 22937 19669 22971 19703
rect 24593 19669 24627 19703
rect 26617 19669 26651 19703
rect 16129 19465 16163 19499
rect 16221 19465 16255 19499
rect 26801 19465 26835 19499
rect 15485 19397 15519 19431
rect 20085 19397 20119 19431
rect 2789 19329 2823 19363
rect 15301 19329 15335 19363
rect 17325 19329 17359 19363
rect 17693 19329 17727 19363
rect 17877 19329 17911 19363
rect 19441 19329 19475 19363
rect 19625 19329 19659 19363
rect 20545 19329 20579 19363
rect 21005 19329 21039 19363
rect 21097 19329 21131 19363
rect 24961 19329 24995 19363
rect 25053 19329 25087 19363
rect 30573 19329 30607 19363
rect 4445 19261 4479 19295
rect 16405 19261 16439 19295
rect 16957 19261 16991 19295
rect 17233 19261 17267 19295
rect 19809 19261 19843 19295
rect 20637 19261 20671 19295
rect 21557 19261 21591 19295
rect 25329 19261 25363 19295
rect 15761 19193 15795 19227
rect 2605 19125 2639 19159
rect 3801 19125 3835 19159
rect 15669 19125 15703 19159
rect 19533 19125 19567 19159
rect 24777 19125 24811 19159
rect 30849 19125 30883 19159
rect 3801 18921 3835 18955
rect 6929 18921 6963 18955
rect 21465 18921 21499 18955
rect 24501 18921 24535 18955
rect 25329 18921 25363 18955
rect 3617 18853 3651 18887
rect 14565 18853 14599 18887
rect 24777 18853 24811 18887
rect 4445 18785 4479 18819
rect 5181 18785 5215 18819
rect 16497 18785 16531 18819
rect 16957 18785 16991 18819
rect 17601 18785 17635 18819
rect 20729 18785 20763 18819
rect 21649 18785 21683 18819
rect 22017 18785 22051 18819
rect 2237 18717 2271 18751
rect 6745 18717 6779 18751
rect 9321 18717 9355 18751
rect 12909 18717 12943 18751
rect 14749 18717 14783 18751
rect 16405 18717 16439 18751
rect 16773 18717 16807 18751
rect 17693 18717 17727 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 21005 18717 21039 18751
rect 25145 18717 25179 18751
rect 2504 18649 2538 18683
rect 4169 18649 4203 18683
rect 4629 18649 4663 18683
rect 15761 18649 15795 18683
rect 17049 18649 17083 18683
rect 21097 18649 21131 18683
rect 21281 18649 21315 18683
rect 24593 18649 24627 18683
rect 24961 18649 24995 18683
rect 4261 18581 4295 18615
rect 9137 18581 9171 18615
rect 12725 18581 12759 18615
rect 20913 18581 20947 18615
rect 21833 18581 21867 18615
rect 3525 18377 3559 18411
rect 3985 18377 4019 18411
rect 4077 18377 4111 18411
rect 6377 18377 6411 18411
rect 6837 18377 6871 18411
rect 10149 18377 10183 18411
rect 15761 18377 15795 18411
rect 18061 18377 18095 18411
rect 23765 18377 23799 18411
rect 25329 18377 25363 18411
rect 8401 18309 8435 18343
rect 9036 18309 9070 18343
rect 12705 18309 12739 18343
rect 16129 18309 16163 18343
rect 18153 18309 18187 18343
rect 23489 18309 23523 18343
rect 24409 18309 24443 18343
rect 1409 18241 1443 18275
rect 2145 18241 2179 18275
rect 2412 18241 2446 18275
rect 4445 18241 4479 18275
rect 4629 18241 4663 18275
rect 4721 18241 4755 18275
rect 4813 18241 4847 18275
rect 6101 18241 6135 18275
rect 6745 18241 6779 18275
rect 7205 18241 7239 18275
rect 8033 18241 8067 18275
rect 10793 18241 10827 18275
rect 12449 18241 12483 18275
rect 15117 18241 15151 18275
rect 15669 18241 15703 18275
rect 16681 18241 16715 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 19257 18241 19291 18275
rect 19441 18241 19475 18275
rect 21281 18241 21315 18275
rect 23305 18241 23339 18275
rect 23949 18241 23983 18275
rect 24041 18241 24075 18275
rect 24685 18241 24719 18275
rect 27077 18241 27111 18275
rect 4261 18173 4295 18207
rect 6929 18173 6963 18207
rect 7849 18173 7883 18207
rect 8769 18173 8803 18207
rect 14289 18173 14323 18207
rect 15301 18173 15335 18207
rect 16221 18173 16255 18207
rect 16405 18173 16439 18207
rect 17325 18173 17359 18207
rect 17601 18173 17635 18207
rect 24225 18173 24259 18207
rect 25053 18173 25087 18207
rect 4997 18105 5031 18139
rect 10241 18105 10275 18139
rect 13829 18105 13863 18139
rect 24850 18105 24884 18139
rect 1593 18037 1627 18071
rect 3617 18037 3651 18071
rect 5917 18037 5951 18071
rect 14841 18037 14875 18071
rect 19441 18037 19475 18071
rect 21373 18037 21407 18071
rect 23121 18037 23155 18071
rect 24041 18037 24075 18071
rect 24317 18037 24351 18071
rect 24961 18037 24995 18071
rect 27169 18037 27203 18071
rect 2513 17833 2547 17867
rect 9321 17833 9355 17867
rect 14105 17833 14139 17867
rect 16037 17833 16071 17867
rect 18889 17833 18923 17867
rect 19349 17833 19383 17867
rect 22569 17833 22603 17867
rect 23949 17833 23983 17867
rect 27813 17833 27847 17867
rect 19993 17765 20027 17799
rect 20637 17765 20671 17799
rect 5457 17697 5491 17731
rect 9781 17697 9815 17731
rect 9873 17697 9907 17731
rect 12449 17697 12483 17731
rect 14565 17697 14599 17731
rect 14749 17697 14783 17731
rect 16129 17697 16163 17731
rect 16773 17697 16807 17731
rect 17785 17697 17819 17731
rect 18981 17697 19015 17731
rect 23397 17697 23431 17731
rect 23489 17697 23523 17731
rect 26065 17697 26099 17731
rect 2697 17629 2731 17663
rect 6929 17629 6963 17663
rect 9689 17629 9723 17663
rect 10977 17629 11011 17663
rect 11345 17629 11379 17663
rect 11713 17629 11747 17663
rect 12173 17629 12207 17663
rect 15853 17629 15887 17663
rect 16313 17629 16347 17663
rect 16635 17629 16669 17663
rect 17969 17629 18003 17663
rect 18521 17629 18555 17663
rect 19073 17629 19107 17663
rect 19441 17629 19475 17663
rect 19549 17639 19583 17673
rect 19809 17629 19843 17663
rect 20085 17629 20119 17663
rect 20361 17629 20395 17663
rect 20453 17629 20487 17663
rect 21189 17629 21223 17663
rect 21373 17629 21407 17663
rect 21925 17629 21959 17663
rect 22201 17629 22235 17663
rect 25513 17629 25547 17663
rect 5724 17561 5758 17595
rect 7174 17561 7208 17595
rect 11437 17561 11471 17595
rect 11529 17561 11563 17595
rect 12694 17561 12728 17595
rect 15669 17561 15703 17595
rect 17325 17561 17359 17595
rect 20269 17561 20303 17595
rect 21741 17561 21775 17595
rect 22753 17561 22787 17595
rect 22937 17561 22971 17595
rect 23581 17561 23615 17595
rect 26341 17561 26375 17595
rect 6837 17493 6871 17527
rect 8309 17493 8343 17527
rect 10425 17493 10459 17527
rect 11161 17493 11195 17527
rect 12357 17493 12391 17527
rect 13829 17493 13863 17527
rect 14473 17493 14507 17527
rect 18705 17493 18739 17527
rect 19625 17493 19659 17527
rect 21373 17493 21407 17527
rect 25697 17493 25731 17527
rect 5917 17289 5951 17323
rect 6837 17289 6871 17323
rect 10149 17289 10183 17323
rect 10701 17289 10735 17323
rect 13001 17289 13035 17323
rect 15209 17289 15243 17323
rect 17141 17289 17175 17323
rect 18429 17289 18463 17323
rect 19533 17289 19567 17323
rect 20821 17289 20855 17323
rect 23397 17289 23431 17323
rect 24409 17289 24443 17323
rect 24869 17289 24903 17323
rect 25237 17289 25271 17323
rect 9036 17221 9070 17255
rect 10609 17221 10643 17255
rect 17049 17221 17083 17255
rect 17693 17221 17727 17255
rect 21833 17221 21867 17255
rect 5733 17153 5767 17187
rect 6745 17153 6779 17187
rect 7205 17153 7239 17187
rect 7849 17153 7883 17187
rect 7941 17153 7975 17187
rect 8034 17153 8068 17187
rect 8217 17153 8251 17187
rect 8309 17153 8343 17187
rect 8447 17153 8481 17187
rect 8769 17153 8803 17187
rect 11529 17153 11563 17187
rect 11713 17153 11747 17187
rect 13369 17153 13403 17187
rect 13829 17153 13863 17187
rect 14381 17153 14415 17187
rect 16497 17153 16531 17187
rect 17969 17153 18003 17187
rect 18245 17153 18279 17187
rect 18521 17153 18555 17187
rect 19165 17153 19199 17187
rect 19257 17153 19291 17187
rect 21005 17153 21039 17187
rect 23581 17153 23615 17187
rect 24041 17153 24075 17187
rect 25329 17153 25363 17187
rect 27169 17153 27203 17187
rect 6929 17085 6963 17119
rect 10885 17085 10919 17119
rect 13461 17085 13495 17119
rect 13645 17085 13679 17119
rect 17233 17085 17267 17119
rect 19073 17085 19107 17119
rect 19349 17085 19383 17119
rect 21097 17085 21131 17119
rect 21189 17085 21223 17119
rect 21281 17085 21315 17119
rect 22201 17085 22235 17119
rect 23765 17085 23799 17119
rect 23949 17085 23983 17119
rect 24593 17085 24627 17119
rect 24777 17085 24811 17119
rect 6377 17017 6411 17051
rect 10241 17017 10275 17051
rect 22109 17017 22143 17051
rect 8585 16949 8619 16983
rect 11529 16949 11563 16983
rect 11897 16949 11931 16983
rect 16681 16949 16715 16983
rect 18061 16949 18095 16983
rect 21998 16949 22032 16983
rect 22477 16949 22511 16983
rect 25513 16949 25547 16983
rect 27077 16949 27111 16983
rect 9137 16745 9171 16779
rect 11161 16745 11195 16779
rect 15853 16745 15887 16779
rect 19441 16745 19475 16779
rect 23673 16745 23707 16779
rect 26138 16745 26172 16779
rect 27629 16745 27663 16779
rect 17417 16677 17451 16711
rect 19625 16677 19659 16711
rect 22753 16677 22787 16711
rect 3065 16609 3099 16643
rect 3249 16609 3283 16643
rect 11805 16609 11839 16643
rect 18429 16609 18463 16643
rect 23305 16609 23339 16643
rect 23489 16609 23523 16643
rect 24409 16609 24443 16643
rect 24685 16609 24719 16643
rect 25881 16609 25915 16643
rect 2513 16541 2547 16575
rect 4353 16541 4387 16575
rect 9321 16541 9355 16575
rect 10517 16541 10551 16575
rect 10665 16541 10699 16575
rect 11023 16541 11057 16575
rect 14105 16541 14139 16575
rect 14473 16541 14507 16575
rect 16037 16541 16071 16575
rect 16313 16541 16347 16575
rect 16681 16541 16715 16575
rect 16773 16541 16807 16575
rect 17509 16541 17543 16575
rect 18797 16541 18831 16575
rect 18981 16541 19015 16575
rect 19717 16541 19751 16575
rect 20729 16541 20763 16575
rect 20913 16541 20947 16575
rect 22937 16541 22971 16575
rect 23029 16541 23063 16575
rect 23213 16541 23247 16575
rect 23397 16541 23431 16575
rect 23857 16541 23891 16575
rect 24777 16541 24811 16575
rect 2973 16473 3007 16507
rect 3801 16473 3835 16507
rect 10793 16473 10827 16507
rect 10885 16473 10919 16507
rect 14289 16473 14323 16507
rect 14381 16473 14415 16507
rect 15485 16473 15519 16507
rect 15669 16473 15703 16507
rect 19257 16473 19291 16507
rect 19809 16473 19843 16507
rect 22753 16473 22787 16507
rect 24225 16473 24259 16507
rect 2329 16405 2363 16439
rect 2605 16405 2639 16439
rect 11253 16405 11287 16439
rect 14657 16405 14691 16439
rect 18797 16405 18831 16439
rect 19457 16405 19491 16439
rect 20821 16405 20855 16439
rect 3341 16201 3375 16235
rect 6837 16201 6871 16235
rect 8677 16201 8711 16235
rect 10241 16201 10275 16235
rect 10609 16201 10643 16235
rect 10701 16201 10735 16235
rect 18245 16201 18279 16235
rect 20913 16201 20947 16235
rect 21373 16201 21407 16235
rect 23305 16201 23339 16235
rect 24685 16201 24719 16235
rect 2228 16133 2262 16167
rect 3893 16133 3927 16167
rect 5181 16133 5215 16167
rect 9014 16133 9048 16167
rect 21281 16133 21315 16167
rect 26341 16133 26375 16167
rect 1685 16065 1719 16099
rect 3801 16065 3835 16099
rect 4261 16065 4295 16099
rect 4997 16065 5031 16099
rect 5273 16065 5307 16099
rect 5365 16065 5399 16099
rect 6745 16065 6779 16099
rect 7205 16065 7239 16099
rect 8493 16065 8527 16099
rect 11989 16065 12023 16099
rect 13001 16065 13035 16099
rect 18153 16065 18187 16099
rect 18337 16065 18371 16099
rect 18797 16065 18831 16099
rect 19257 16065 19291 16099
rect 19533 16065 19567 16099
rect 19809 16065 19843 16099
rect 20085 16065 20119 16099
rect 23213 16065 23247 16099
rect 23397 16065 23431 16099
rect 23489 16065 23523 16099
rect 23857 16065 23891 16099
rect 24317 16065 24351 16099
rect 26157 16065 26191 16099
rect 26433 16065 26467 16099
rect 26525 16065 26559 16099
rect 1961 15997 1995 16031
rect 3985 15997 4019 16031
rect 4813 15997 4847 16031
rect 6929 15997 6963 16031
rect 7849 15997 7883 16031
rect 8769 15997 8803 16031
rect 10793 15997 10827 16031
rect 13277 15997 13311 16031
rect 18521 15997 18555 16031
rect 19901 15997 19935 16031
rect 21465 15997 21499 16031
rect 24225 15997 24259 16031
rect 3433 15929 3467 15963
rect 5549 15929 5583 15963
rect 10149 15929 10183 15963
rect 1869 15861 1903 15895
rect 6377 15861 6411 15895
rect 12173 15861 12207 15895
rect 12817 15861 12851 15895
rect 13185 15861 13219 15895
rect 26709 15861 26743 15895
rect 3433 15657 3467 15691
rect 8309 15657 8343 15691
rect 13645 15657 13679 15691
rect 19441 15657 19475 15691
rect 23029 15657 23063 15691
rect 28549 15657 28583 15691
rect 17969 15589 18003 15623
rect 11253 15521 11287 15555
rect 12265 15521 12299 15555
rect 14657 15521 14691 15555
rect 18521 15521 18555 15555
rect 18613 15521 18647 15555
rect 28365 15521 28399 15555
rect 29193 15521 29227 15555
rect 2053 15453 2087 15487
rect 5181 15453 5215 15487
rect 5457 15453 5491 15487
rect 6929 15453 6963 15487
rect 9229 15453 9263 15487
rect 12081 15453 12115 15487
rect 12521 15453 12555 15487
rect 15853 15453 15887 15487
rect 17693 15453 17727 15487
rect 17785 15453 17819 15487
rect 21005 15453 21039 15487
rect 21281 15453 21315 15487
rect 26065 15453 26099 15487
rect 27721 15453 27755 15487
rect 19487 15419 19521 15453
rect 2298 15385 2332 15419
rect 5724 15385 5758 15419
rect 7174 15385 7208 15419
rect 9496 15385 9530 15419
rect 17969 15385 18003 15419
rect 19257 15385 19291 15419
rect 21557 15385 21591 15419
rect 26893 15385 26927 15419
rect 5365 15317 5399 15351
rect 6837 15317 6871 15351
rect 10609 15317 10643 15351
rect 10701 15317 10735 15351
rect 11069 15317 11103 15351
rect 11161 15317 11195 15351
rect 11529 15317 11563 15351
rect 14105 15317 14139 15351
rect 15301 15317 15335 15351
rect 18061 15317 18095 15351
rect 18429 15317 18463 15351
rect 19625 15317 19659 15351
rect 21189 15317 21223 15351
rect 26709 15317 26743 15351
rect 27813 15317 27847 15351
rect 5825 15113 5859 15147
rect 6837 15113 6871 15147
rect 9597 15113 9631 15147
rect 12817 15113 12851 15147
rect 13185 15113 13219 15147
rect 13277 15113 13311 15147
rect 14933 15113 14967 15147
rect 15025 15113 15059 15147
rect 16497 15113 16531 15147
rect 21925 15113 21959 15147
rect 25513 15113 25547 15147
rect 26341 15113 26375 15147
rect 26801 15113 26835 15147
rect 29193 15113 29227 15147
rect 8217 15045 8251 15079
rect 27721 15045 27755 15079
rect 29377 15045 29411 15079
rect 6009 14977 6043 15011
rect 6745 14977 6779 15011
rect 7205 14977 7239 15011
rect 7757 14977 7791 15011
rect 7941 14977 7975 15011
rect 8089 14977 8123 15011
rect 8309 14977 8343 15011
rect 8447 14977 8481 15011
rect 9781 14977 9815 15011
rect 15393 14977 15427 15011
rect 15541 14977 15575 15011
rect 15669 14977 15703 15011
rect 15761 14977 15795 15011
rect 15858 14977 15892 15011
rect 16129 14977 16163 15011
rect 17693 14977 17727 15011
rect 18613 14977 18647 15011
rect 18797 14977 18831 15011
rect 18889 14977 18923 15011
rect 20545 14977 20579 15011
rect 21281 14977 21315 15011
rect 22017 14977 22051 15011
rect 25697 14977 25731 15011
rect 26433 14977 26467 15011
rect 26985 14977 27019 15011
rect 29469 14977 29503 15011
rect 6929 14909 6963 14943
rect 12449 14909 12483 14943
rect 13461 14909 13495 14943
rect 14197 14909 14231 14943
rect 15117 14909 15151 14943
rect 16221 14909 16255 14943
rect 18429 14909 18463 14943
rect 25973 14909 26007 14943
rect 26249 14909 26283 14943
rect 27445 14909 27479 14943
rect 6377 14841 6411 14875
rect 8585 14841 8619 14875
rect 16037 14841 16071 14875
rect 11897 14773 11931 14807
rect 13645 14773 13679 14807
rect 14565 14773 14599 14807
rect 16129 14773 16163 14807
rect 17509 14773 17543 14807
rect 19073 14773 19107 14807
rect 20637 14773 20671 14807
rect 25881 14773 25915 14807
rect 27169 14773 27203 14807
rect 15577 14569 15611 14603
rect 18613 14569 18647 14603
rect 26341 14569 26375 14603
rect 13921 14501 13955 14535
rect 11621 14433 11655 14467
rect 11897 14433 11931 14467
rect 17141 14433 17175 14467
rect 13645 14365 13679 14399
rect 13737 14365 13771 14399
rect 14197 14365 14231 14399
rect 16865 14365 16899 14399
rect 27721 14365 27755 14399
rect 13553 14297 13587 14331
rect 14442 14297 14476 14331
rect 27454 14297 27488 14331
rect 13369 14229 13403 14263
rect 3065 14025 3099 14059
rect 8861 14025 8895 14059
rect 11897 14025 11931 14059
rect 14289 14025 14323 14059
rect 15761 14025 15795 14059
rect 17877 14025 17911 14059
rect 24777 14025 24811 14059
rect 12173 13957 12207 13991
rect 12265 13957 12299 13991
rect 14626 13957 14660 13991
rect 2513 13889 2547 13923
rect 2973 13889 3007 13923
rect 3433 13889 3467 13923
rect 8677 13889 8711 13923
rect 12081 13889 12115 13923
rect 12449 13889 12483 13923
rect 14105 13889 14139 13923
rect 16405 13889 16439 13923
rect 17785 13889 17819 13923
rect 24409 13889 24443 13923
rect 3157 13821 3191 13855
rect 3985 13821 4019 13855
rect 9689 13821 9723 13855
rect 14381 13821 14415 13855
rect 24501 13821 24535 13855
rect 2329 13685 2363 13719
rect 2605 13685 2639 13719
rect 9137 13685 9171 13719
rect 15853 13685 15887 13719
rect 24409 13685 24443 13719
rect 3801 13481 3835 13515
rect 8769 13481 8803 13515
rect 14841 13481 14875 13515
rect 30573 13481 30607 13515
rect 3341 13413 3375 13447
rect 4261 13345 4295 13379
rect 4445 13345 4479 13379
rect 6561 13345 6595 13379
rect 9413 13345 9447 13379
rect 9505 13345 9539 13379
rect 15393 13345 15427 13379
rect 22753 13345 22787 13379
rect 24961 13345 24995 13379
rect 1685 13277 1719 13311
rect 1961 13277 1995 13311
rect 5181 13277 5215 13311
rect 5549 13277 5583 13311
rect 5825 13277 5859 13311
rect 5973 13277 6007 13311
rect 6331 13277 6365 13311
rect 7389 13277 7423 13311
rect 9321 13277 9355 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 11069 13277 11103 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 23489 13277 23523 13311
rect 25789 13277 25823 13311
rect 2206 13209 2240 13243
rect 4169 13209 4203 13243
rect 4629 13209 4663 13243
rect 6101 13209 6135 13243
rect 6193 13209 6227 13243
rect 7656 13209 7690 13243
rect 10885 13209 10919 13243
rect 30849 13209 30883 13243
rect 1869 13141 1903 13175
rect 5365 13141 5399 13175
rect 6469 13141 6503 13175
rect 7205 13141 7239 13175
rect 8953 13141 8987 13175
rect 9965 13141 9999 13175
rect 11253 13141 11287 13175
rect 22109 13141 22143 13175
rect 22477 13141 22511 13175
rect 22569 13141 22603 13175
rect 22937 13141 22971 13175
rect 24409 13141 24443 13175
rect 24777 13141 24811 13175
rect 24869 13141 24903 13175
rect 25237 13141 25271 13175
rect 3341 12937 3375 12971
rect 4169 12937 4203 12971
rect 6193 12937 6227 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 9413 12937 9447 12971
rect 9505 12937 9539 12971
rect 19441 12937 19475 12971
rect 21373 12937 21407 12971
rect 21649 12937 21683 12971
rect 23213 12937 23247 12971
rect 23765 12937 23799 12971
rect 25237 12937 25271 12971
rect 3893 12869 3927 12903
rect 6837 12869 6871 12903
rect 7941 12869 7975 12903
rect 8769 12869 8803 12903
rect 11253 12869 11287 12903
rect 21005 12869 21039 12903
rect 22078 12869 22112 12903
rect 24102 12869 24136 12903
rect 25697 12869 25731 12903
rect 1961 12801 1995 12835
rect 2228 12801 2262 12835
rect 3617 12801 3651 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 4813 12801 4847 12835
rect 5080 12801 5114 12835
rect 10425 12801 10459 12835
rect 17049 12801 17083 12835
rect 19073 12801 19107 12835
rect 19533 12801 19567 12835
rect 19993 12801 20027 12835
rect 20729 12801 20763 12835
rect 20822 12801 20856 12835
rect 21097 12801 21131 12835
rect 21194 12801 21228 12835
rect 21465 12801 21499 12835
rect 21833 12801 21867 12835
rect 23305 12801 23339 12835
rect 23581 12801 23615 12835
rect 25789 12801 25823 12835
rect 26157 12801 26191 12835
rect 28641 12801 28675 12835
rect 6929 12733 6963 12767
rect 9597 12733 9631 12767
rect 13185 12733 13219 12767
rect 17141 12733 17175 12767
rect 17325 12733 17359 12767
rect 18153 12733 18187 12767
rect 19349 12733 19383 12767
rect 20637 12733 20671 12767
rect 23857 12733 23891 12767
rect 25881 12733 25915 12767
rect 26709 12733 26743 12767
rect 28089 12733 28123 12767
rect 9045 12597 9079 12631
rect 13737 12597 13771 12631
rect 16681 12597 16715 12631
rect 17601 12597 17635 12631
rect 18429 12597 18463 12631
rect 19901 12597 19935 12631
rect 23489 12597 23523 12631
rect 25329 12597 25363 12631
rect 27445 12597 27479 12631
rect 28549 12597 28583 12631
rect 8217 12393 8251 12427
rect 10333 12393 10367 12427
rect 11437 12393 11471 12427
rect 17509 12393 17543 12427
rect 19073 12393 19107 12427
rect 20637 12393 20671 12427
rect 24225 12393 24259 12427
rect 25789 12393 25823 12427
rect 29101 12393 29135 12427
rect 6469 12325 6503 12359
rect 11253 12325 11287 12359
rect 11713 12325 11747 12359
rect 5089 12257 5123 12291
rect 7021 12257 7055 12291
rect 7113 12257 7147 12291
rect 7941 12257 7975 12291
rect 11437 12257 11471 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 17325 12257 17359 12291
rect 18429 12257 18463 12291
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 8953 12189 8987 12223
rect 10609 12189 10643 12223
rect 10702 12189 10736 12223
rect 10977 12189 11011 12223
rect 11074 12189 11108 12223
rect 11345 12189 11379 12223
rect 12265 12189 12299 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 17049 12189 17083 12223
rect 18061 12189 18095 12223
rect 18705 12189 18739 12223
rect 19257 12189 19291 12223
rect 20913 12189 20947 12223
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 22957 12189 22991 12223
rect 23305 12189 23339 12223
rect 23581 12189 23615 12223
rect 23729 12189 23763 12223
rect 23949 12189 23983 12223
rect 24087 12189 24121 12223
rect 24409 12189 24443 12223
rect 26433 12189 26467 12223
rect 26525 12189 26559 12223
rect 26709 12189 26743 12223
rect 27353 12189 27387 12223
rect 5356 12121 5390 12155
rect 9198 12121 9232 12155
rect 10885 12121 10919 12155
rect 12357 12121 12391 12155
rect 19524 12121 19558 12155
rect 21732 12121 21766 12155
rect 23121 12121 23155 12155
rect 23213 12121 23247 12155
rect 23857 12121 23891 12155
rect 24654 12121 24688 12155
rect 27629 12121 27663 12155
rect 6561 12053 6595 12087
rect 6929 12053 6963 12087
rect 7389 12053 7423 12087
rect 8769 12053 8803 12087
rect 12081 12053 12115 12087
rect 13461 12053 13495 12087
rect 13829 12053 13863 12087
rect 16681 12053 16715 12087
rect 17141 12053 17175 12087
rect 18613 12053 18647 12087
rect 20729 12053 20763 12087
rect 21005 12053 21039 12087
rect 22845 12053 22879 12087
rect 23489 12053 23523 12087
rect 26893 12053 26927 12087
rect 5549 11849 5583 11883
rect 8861 11849 8895 11883
rect 14197 11849 14231 11883
rect 15393 11849 15427 11883
rect 18061 11849 18095 11883
rect 18981 11849 19015 11883
rect 21649 11849 21683 11883
rect 26065 11849 26099 11883
rect 26525 11849 26559 11883
rect 28365 11849 28399 11883
rect 22661 11781 22695 11815
rect 1409 11713 1443 11747
rect 1777 11713 1811 11747
rect 3985 11713 4019 11747
rect 5733 11713 5767 11747
rect 8585 11713 8619 11747
rect 9229 11713 9263 11747
rect 9689 11713 9723 11747
rect 9956 11713 9990 11747
rect 11345 11713 11379 11747
rect 12081 11713 12115 11747
rect 13849 11713 13883 11747
rect 14105 11713 14139 11747
rect 14749 11713 14783 11747
rect 15025 11713 15059 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 16221 11713 16255 11747
rect 16313 11713 16347 11747
rect 16681 11713 16715 11747
rect 16937 11713 16971 11747
rect 18153 11713 18187 11747
rect 18337 11713 18371 11747
rect 18429 11713 18463 11747
rect 18521 11713 18555 11747
rect 20105 11713 20139 11747
rect 20361 11713 20395 11747
rect 21465 11713 21499 11747
rect 21833 11713 21867 11747
rect 23397 11713 23431 11747
rect 25789 11713 25823 11747
rect 26433 11713 26467 11747
rect 27241 11713 27275 11747
rect 9321 11645 9355 11679
rect 9505 11645 9539 11679
rect 14933 11645 14967 11679
rect 26709 11645 26743 11679
rect 26985 11645 27019 11679
rect 29101 11645 29135 11679
rect 11161 11577 11195 11611
rect 15485 11577 15519 11611
rect 16497 11577 16531 11611
rect 25973 11577 26007 11611
rect 3801 11509 3835 11543
rect 8769 11509 8803 11543
rect 11069 11509 11103 11543
rect 12633 11509 12667 11543
rect 12725 11509 12759 11543
rect 16037 11509 16071 11543
rect 18705 11509 18739 11543
rect 22845 11509 22879 11543
rect 28457 11509 28491 11543
rect 10333 11305 10367 11339
rect 11161 11305 11195 11339
rect 13921 11305 13955 11339
rect 17325 11305 17359 11339
rect 21833 11305 21867 11339
rect 27261 11305 27295 11339
rect 3617 11237 3651 11271
rect 2237 11169 2271 11203
rect 4537 11169 4571 11203
rect 8953 11169 8987 11203
rect 10609 11169 10643 11203
rect 11805 11169 11839 11203
rect 12449 11169 12483 11203
rect 19441 11169 19475 11203
rect 22477 11169 22511 11203
rect 4997 11101 5031 11135
rect 9209 11101 9243 11135
rect 10793 11101 10827 11135
rect 12173 11101 12207 11135
rect 14289 11101 14323 11135
rect 15945 11101 15979 11135
rect 22201 11101 22235 11135
rect 26709 11101 26743 11135
rect 26985 11101 27019 11135
rect 27077 11101 27111 11135
rect 2504 11033 2538 11067
rect 3985 11033 4019 11067
rect 10701 11033 10735 11067
rect 11253 11033 11287 11067
rect 14197 11033 14231 11067
rect 16190 11033 16224 11067
rect 20177 11033 20211 11067
rect 22293 11033 22327 11067
rect 26893 11033 26927 11067
rect 5641 10965 5675 10999
rect 2973 10761 3007 10795
rect 4721 10761 4755 10795
rect 4813 10761 4847 10795
rect 5181 10761 5215 10795
rect 9873 10761 9907 10795
rect 24777 10761 24811 10795
rect 3608 10693 3642 10727
rect 5273 10693 5307 10727
rect 3157 10625 3191 10659
rect 10517 10625 10551 10659
rect 24409 10625 24443 10659
rect 3341 10557 3375 10591
rect 5365 10557 5399 10591
rect 24501 10557 24535 10591
rect 24409 10421 24443 10455
rect 3801 10217 3835 10251
rect 4261 10081 4295 10115
rect 4353 10081 4387 10115
rect 19993 10081 20027 10115
rect 25973 10081 26007 10115
rect 4169 10013 4203 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 5089 10013 5123 10047
rect 5181 10013 5215 10047
rect 7757 10013 7791 10047
rect 10425 10013 10459 10047
rect 18061 10013 18095 10047
rect 20821 10013 20855 10047
rect 22937 10013 22971 10047
rect 23305 10013 23339 10047
rect 25237 10013 25271 10047
rect 19809 9945 19843 9979
rect 20269 9945 20303 9979
rect 23121 9945 23155 9979
rect 23213 9945 23247 9979
rect 5365 9877 5399 9911
rect 7205 9877 7239 9911
rect 9873 9877 9907 9911
rect 17417 9877 17451 9911
rect 19441 9877 19475 9911
rect 19901 9877 19935 9911
rect 23489 9877 23523 9911
rect 24685 9877 24719 9911
rect 25421 9877 25455 9911
rect 6929 9673 6963 9707
rect 9689 9673 9723 9707
rect 17141 9673 17175 9707
rect 21373 9673 21407 9707
rect 24409 9673 24443 9707
rect 24777 9673 24811 9707
rect 25605 9673 25639 9707
rect 7021 9605 7055 9639
rect 7665 9605 7699 9639
rect 9229 9605 9263 9639
rect 10425 9605 10459 9639
rect 22477 9605 22511 9639
rect 24133 9605 24167 9639
rect 2513 9537 2547 9571
rect 2973 9537 3007 9571
rect 3433 9537 3467 9571
rect 7389 9537 7423 9571
rect 7537 9537 7571 9571
rect 7757 9537 7791 9571
rect 7854 9537 7888 9571
rect 11253 9537 11287 9571
rect 12265 9537 12299 9571
rect 15945 9537 15979 9571
rect 18061 9537 18095 9571
rect 18521 9537 18555 9571
rect 19513 9537 19547 9571
rect 20729 9537 20763 9571
rect 20822 9537 20856 9571
rect 21005 9537 21039 9571
rect 21097 9537 21131 9571
rect 21194 9537 21228 9571
rect 22385 9537 22419 9571
rect 22845 9537 22879 9571
rect 23397 9537 23431 9571
rect 23765 9537 23799 9571
rect 23913 9537 23947 9571
rect 24041 9537 24075 9571
rect 24230 9537 24264 9571
rect 24869 9537 24903 9571
rect 25697 9537 25731 9571
rect 26157 9537 26191 9571
rect 3065 9469 3099 9503
rect 3157 9469 3191 9503
rect 4077 9469 4111 9503
rect 7113 9469 7147 9503
rect 8401 9469 8435 9503
rect 9781 9469 9815 9503
rect 9965 9469 9999 9503
rect 12081 9469 12115 9503
rect 12357 9469 12391 9503
rect 17233 9469 17267 9503
rect 17325 9469 17359 9503
rect 18153 9469 18187 9503
rect 18337 9469 18371 9503
rect 19073 9469 19107 9503
rect 19257 9469 19291 9503
rect 22661 9469 22695 9503
rect 24593 9469 24627 9503
rect 25421 9469 25455 9503
rect 2605 9401 2639 9435
rect 16773 9401 16807 9435
rect 20637 9401 20671 9435
rect 26341 9401 26375 9435
rect 2329 9333 2363 9367
rect 6561 9333 6595 9367
rect 8033 9333 8067 9367
rect 9321 9333 9355 9367
rect 11529 9333 11563 9367
rect 12265 9333 12299 9367
rect 12633 9333 12667 9367
rect 16129 9333 16163 9367
rect 17693 9333 17727 9367
rect 22017 9333 22051 9367
rect 25237 9333 25271 9367
rect 26065 9333 26099 9367
rect 7389 9129 7423 9163
rect 12265 9129 12299 9163
rect 19073 9129 19107 9163
rect 20637 9129 20671 9163
rect 23121 9129 23155 9163
rect 24409 9129 24443 9163
rect 3341 9061 3375 9095
rect 5917 9061 5951 9095
rect 10885 9061 10919 9095
rect 23949 9061 23983 9095
rect 25881 9061 25915 9095
rect 6009 8993 6043 9027
rect 8033 8993 8067 9027
rect 12909 8993 12943 9027
rect 19257 8993 19291 9027
rect 23305 8993 23339 9027
rect 1961 8925 1995 8959
rect 4629 8925 4663 8959
rect 5457 8925 5491 8959
rect 5733 8925 5767 8959
rect 6265 8925 6299 8959
rect 7941 8925 7975 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9505 8925 9539 8959
rect 10977 8925 11011 8959
rect 11161 8925 11195 8959
rect 11345 8925 11379 8959
rect 11621 8925 11655 8959
rect 11769 8925 11803 8959
rect 12086 8925 12120 8959
rect 12725 8925 12759 8959
rect 13737 8925 13771 8959
rect 16037 8925 16071 8959
rect 16221 8925 16255 8959
rect 17969 8925 18003 8959
rect 18797 8925 18831 8959
rect 18889 8925 18923 8959
rect 20821 8925 20855 8959
rect 21741 8925 21775 8959
rect 24225 8925 24259 8959
rect 25533 8925 25567 8959
rect 25789 8925 25823 8959
rect 26065 8925 26099 8959
rect 26341 8925 26375 8959
rect 2228 8857 2262 8891
rect 9750 8857 9784 8891
rect 11253 8857 11287 8891
rect 11897 8857 11931 8891
rect 11989 8857 12023 8891
rect 16466 8857 16500 8891
rect 19524 8857 19558 8891
rect 21649 8857 21683 8891
rect 21986 8857 22020 8891
rect 23581 8857 23615 8891
rect 4077 8789 4111 8823
rect 5641 8789 5675 8823
rect 7481 8789 7515 8823
rect 7849 8789 7883 8823
rect 8953 8789 8987 8823
rect 9413 8789 9447 8823
rect 11529 8789 11563 8823
rect 12357 8789 12391 8823
rect 12817 8789 12851 8823
rect 13185 8789 13219 8823
rect 15485 8789 15519 8823
rect 17601 8789 17635 8823
rect 23489 8789 23523 8823
rect 24041 8789 24075 8823
rect 26157 8789 26191 8823
rect 3801 8585 3835 8619
rect 4261 8585 4295 8619
rect 7757 8585 7791 8619
rect 7849 8585 7883 8619
rect 10057 8585 10091 8619
rect 10517 8585 10551 8619
rect 11897 8585 11931 8619
rect 13369 8585 13403 8619
rect 15301 8585 15335 8619
rect 15669 8585 15703 8619
rect 16497 8585 16531 8619
rect 18061 8585 18095 8619
rect 19625 8585 19659 8619
rect 20913 8585 20947 8619
rect 21649 8585 21683 8619
rect 23581 8585 23615 8619
rect 24593 8585 24627 8619
rect 4997 8517 5031 8551
rect 12256 8517 12290 8551
rect 16926 8517 16960 8551
rect 18705 8517 18739 8551
rect 18797 8517 18831 8551
rect 2421 8449 2455 8483
rect 2688 8449 2722 8483
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 5089 8449 5123 8483
rect 6377 8449 6411 8483
rect 6633 8449 6667 8483
rect 8401 8449 8435 8483
rect 8585 8449 8619 8483
rect 8852 8449 8886 8483
rect 10425 8449 10459 8483
rect 11161 8449 11195 8483
rect 11713 8449 11747 8483
rect 11989 8449 12023 8483
rect 13829 8449 13863 8483
rect 13921 8449 13955 8483
rect 14289 8449 14323 8483
rect 14841 8449 14875 8483
rect 15209 8449 15243 8483
rect 15761 8449 15795 8483
rect 16313 8449 16347 8483
rect 16681 8449 16715 8483
rect 18521 8449 18555 8483
rect 18889 8449 18923 8483
rect 19717 8449 19751 8483
rect 20177 8449 20211 8483
rect 20821 8449 20855 8483
rect 21097 8449 21131 8483
rect 21465 8449 21499 8483
rect 22376 8449 22410 8483
rect 25717 8449 25751 8483
rect 25973 8449 26007 8483
rect 4353 8381 4387 8415
rect 4445 8381 4479 8415
rect 10609 8381 10643 8415
rect 14105 8381 14139 8415
rect 15945 8381 15979 8415
rect 19533 8381 19567 8415
rect 22109 8381 22143 8415
rect 24133 8381 24167 8415
rect 5273 8313 5307 8347
rect 9965 8313 9999 8347
rect 13461 8313 13495 8347
rect 19073 8313 19107 8347
rect 20085 8313 20119 8347
rect 23489 8313 23523 8347
rect 3893 8245 3927 8279
rect 11345 8245 11379 8279
rect 15025 8245 15059 8279
rect 2697 8041 2731 8075
rect 7205 8041 7239 8075
rect 12909 8041 12943 8075
rect 30757 8041 30791 8075
rect 16129 7973 16163 8007
rect 18337 7973 18371 8007
rect 16865 7905 16899 7939
rect 2881 7837 2915 7871
rect 6929 7837 6963 7871
rect 11529 7837 11563 7871
rect 14473 7837 14507 7871
rect 14749 7837 14783 7871
rect 15016 7837 15050 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 18061 7837 18095 7871
rect 18153 7837 18187 7871
rect 30941 7837 30975 7871
rect 11774 7769 11808 7803
rect 16589 7769 16623 7803
rect 17049 7769 17083 7803
rect 17969 7769 18003 7803
rect 14657 7701 14691 7735
rect 16221 7701 16255 7735
rect 16681 7701 16715 7735
rect 16313 7497 16347 7531
rect 15178 7429 15212 7463
rect 14933 7361 14967 7395
rect 25145 6953 25179 6987
rect 19073 6885 19107 6919
rect 6929 6817 6963 6851
rect 7941 6817 7975 6851
rect 19809 6817 19843 6851
rect 21833 6817 21867 6851
rect 6101 6749 6135 6783
rect 8033 6749 8067 6783
rect 8126 6749 8160 6783
rect 8309 6749 8343 6783
rect 8401 6749 8435 6783
rect 8498 6749 8532 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 18429 6749 18463 6783
rect 18577 6749 18611 6783
rect 18705 6749 18739 6783
rect 18935 6749 18969 6783
rect 20729 6749 20763 6783
rect 21097 6749 21131 6783
rect 21649 6749 21683 6783
rect 22201 6749 22235 6783
rect 22569 6749 22603 6783
rect 24409 6749 24443 6783
rect 24502 6749 24536 6783
rect 24685 6749 24719 6783
rect 24874 6749 24908 6783
rect 25145 6749 25179 6783
rect 25237 6749 25271 6783
rect 6745 6681 6779 6715
rect 7297 6681 7331 6715
rect 10885 6681 10919 6715
rect 18797 6681 18831 6715
rect 19625 6681 19659 6715
rect 20085 6681 20119 6715
rect 22385 6681 22419 6715
rect 22477 6681 22511 6715
rect 24777 6681 24811 6715
rect 6285 6613 6319 6647
rect 6377 6613 6411 6647
rect 6837 6613 6871 6647
rect 8677 6613 8711 6647
rect 9965 6613 9999 6647
rect 11253 6613 11287 6647
rect 19257 6613 19291 6647
rect 19717 6613 19751 6647
rect 20913 6613 20947 6647
rect 21189 6613 21223 6647
rect 21557 6613 21591 6647
rect 22753 6613 22787 6647
rect 25053 6613 25087 6647
rect 25513 6613 25547 6647
rect 5457 6409 5491 6443
rect 5917 6409 5951 6443
rect 7757 6409 7791 6443
rect 8033 6409 8067 6443
rect 9689 6409 9723 6443
rect 10149 6409 10183 6443
rect 14105 6409 14139 6443
rect 20821 6409 20855 6443
rect 21925 6409 21959 6443
rect 23765 6409 23799 6443
rect 24593 6409 24627 6443
rect 23673 6341 23707 6375
rect 25053 6341 25087 6375
rect 5181 6273 5215 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6633 6273 6667 6307
rect 7849 6273 7883 6307
rect 8309 6273 8343 6307
rect 8576 6273 8610 6307
rect 11529 6273 11563 6307
rect 13461 6273 13495 6307
rect 14197 6273 14231 6307
rect 14565 6273 14599 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 18236 6273 18270 6307
rect 19441 6273 19475 6307
rect 19697 6273 19731 6307
rect 23213 6273 23247 6307
rect 24685 6273 24719 6307
rect 25789 6273 25823 6307
rect 26341 6273 26375 6307
rect 6101 6205 6135 6239
rect 10241 6205 10275 6239
rect 10333 6205 10367 6239
rect 11161 6205 11195 6239
rect 11621 6205 11655 6239
rect 14289 6205 14323 6239
rect 15209 6205 15243 6239
rect 21465 6205 21499 6239
rect 22477 6205 22511 6239
rect 23581 6205 23615 6239
rect 24777 6205 24811 6239
rect 25605 6205 25639 6239
rect 13737 6137 13771 6171
rect 20913 6137 20947 6171
rect 5365 6069 5399 6103
rect 9781 6069 9815 6103
rect 10609 6069 10643 6103
rect 11529 6069 11563 6103
rect 11897 6069 11931 6103
rect 13645 6069 13679 6103
rect 17877 6069 17911 6103
rect 19349 6069 19383 6103
rect 22661 6069 22695 6103
rect 24133 6069 24167 6103
rect 24225 6069 24259 6103
rect 7113 5865 7147 5899
rect 8953 5865 8987 5899
rect 11989 5865 12023 5899
rect 15485 5865 15519 5899
rect 18337 5865 18371 5899
rect 22109 5865 22143 5899
rect 23581 5865 23615 5899
rect 25789 5865 25823 5899
rect 7021 5797 7055 5831
rect 25881 5797 25915 5831
rect 5641 5729 5675 5763
rect 7757 5729 7791 5763
rect 10149 5729 10183 5763
rect 10333 5729 10367 5763
rect 11161 5729 11195 5763
rect 19901 5729 19935 5763
rect 26525 5729 26559 5763
rect 1409 5661 1443 5695
rect 5897 5661 5931 5695
rect 9137 5661 9171 5695
rect 11345 5661 11379 5695
rect 11438 5661 11472 5695
rect 11621 5661 11655 5695
rect 11851 5661 11885 5695
rect 14105 5661 14139 5695
rect 18521 5661 18555 5695
rect 19625 5661 19659 5695
rect 20729 5661 20763 5695
rect 20996 5661 21030 5695
rect 22201 5661 22235 5695
rect 23857 5661 23891 5695
rect 23949 5661 23983 5695
rect 24409 5661 24443 5695
rect 26249 5661 26283 5695
rect 27261 5661 27295 5695
rect 10057 5593 10091 5627
rect 10885 5593 10919 5627
rect 11713 5593 11747 5627
rect 14350 5593 14384 5627
rect 22446 5593 22480 5627
rect 24654 5593 24688 5627
rect 1593 5525 1627 5559
rect 9689 5525 9723 5559
rect 10517 5525 10551 5559
rect 10977 5525 11011 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 23673 5525 23707 5559
rect 24133 5525 24167 5559
rect 26341 5525 26375 5559
rect 26709 5525 26743 5559
rect 10609 5321 10643 5355
rect 11529 5321 11563 5355
rect 21833 5321 21867 5355
rect 22201 5321 22235 5355
rect 22293 5321 22327 5355
rect 24317 5321 24351 5355
rect 25329 5321 25363 5355
rect 12909 5253 12943 5287
rect 13001 5253 13035 5287
rect 13369 5253 13403 5287
rect 25666 5253 25700 5287
rect 9229 5185 9263 5219
rect 9485 5185 9519 5219
rect 12633 5185 12667 5219
rect 12725 5185 12759 5219
rect 13093 5185 13127 5219
rect 15025 5185 15059 5219
rect 15301 5185 15335 5219
rect 21189 5185 21223 5219
rect 22937 5185 22971 5219
rect 23204 5185 23238 5219
rect 25145 5185 25179 5219
rect 25421 5185 25455 5219
rect 27261 5185 27295 5219
rect 12081 5117 12115 5151
rect 13921 5117 13955 5151
rect 14657 5117 14691 5151
rect 22477 5117 22511 5151
rect 26985 5117 27019 5151
rect 14841 5049 14875 5083
rect 15209 5049 15243 5083
rect 21373 5049 21407 5083
rect 26801 5049 26835 5083
rect 12449 4981 12483 5015
rect 13277 4981 13311 5015
rect 14105 4981 14139 5015
rect 27077 4981 27111 5015
rect 27445 4981 27479 5015
rect 9505 4777 9539 4811
rect 13093 4777 13127 4811
rect 15117 4777 15151 4811
rect 17785 4777 17819 4811
rect 9413 4709 9447 4743
rect 10057 4709 10091 4743
rect 12265 4709 12299 4743
rect 26617 4709 26651 4743
rect 10701 4641 10735 4675
rect 12357 4641 12391 4675
rect 13553 4641 13587 4675
rect 13737 4641 13771 4675
rect 14289 4641 14323 4675
rect 16589 4641 16623 4675
rect 18153 4641 18187 4675
rect 26985 4641 27019 4675
rect 9229 4573 9263 4607
rect 9689 4573 9723 4607
rect 9965 4573 9999 4607
rect 10425 4573 10459 4607
rect 11713 4573 11747 4607
rect 11897 4573 11931 4607
rect 12081 4573 12115 4607
rect 13461 4573 13495 4607
rect 15025 4573 15059 4607
rect 15301 4573 15335 4607
rect 15485 4573 15519 4607
rect 15761 4573 15795 4607
rect 16405 4573 16439 4607
rect 17049 4573 17083 4607
rect 17417 4573 17451 4607
rect 17693 4573 17727 4607
rect 17969 4573 18003 4607
rect 26065 4573 26099 4607
rect 26249 4573 26283 4607
rect 26433 4573 26467 4607
rect 28365 4573 28399 4607
rect 11989 4505 12023 4539
rect 17233 4505 17267 4539
rect 17325 4505 17359 4539
rect 26341 4505 26375 4539
rect 27721 4505 27755 4539
rect 9781 4437 9815 4471
rect 10517 4437 10551 4471
rect 13001 4437 13035 4471
rect 14933 4437 14967 4471
rect 15945 4437 15979 4471
rect 16037 4437 16071 4471
rect 16497 4437 16531 4471
rect 17601 4437 17635 4471
rect 27629 4437 27663 4471
rect 15301 4233 15335 4267
rect 16865 4233 16899 4267
rect 18429 4233 18463 4267
rect 14841 4165 14875 4199
rect 9321 4097 9355 4131
rect 9588 4097 9622 4131
rect 11897 4097 11931 4131
rect 12164 4097 12198 4131
rect 15117 4097 15151 4131
rect 15393 4097 15427 4131
rect 17509 4097 17543 4131
rect 18245 4097 18279 4131
rect 26985 4097 27019 4131
rect 13369 4029 13403 4063
rect 19073 4029 19107 4063
rect 27261 4029 27295 4063
rect 10701 3961 10735 3995
rect 13277 3893 13311 3927
rect 17693 3893 17727 3927
rect 28733 3893 28767 3927
rect 10885 3689 10919 3723
rect 14105 3689 14139 3723
rect 17141 3689 17175 3723
rect 27261 3689 27295 3723
rect 10793 3621 10827 3655
rect 11529 3553 11563 3587
rect 12173 3553 12207 3587
rect 12449 3553 12483 3587
rect 13921 3553 13955 3587
rect 14657 3553 14691 3587
rect 15761 3553 15795 3587
rect 17601 3553 17635 3587
rect 19349 3553 19383 3587
rect 9413 3485 9447 3519
rect 15025 3485 15059 3519
rect 16028 3485 16062 3519
rect 17325 3485 17359 3519
rect 19441 3485 19475 3519
rect 27169 3485 27203 3519
rect 9680 3417 9714 3451
rect 14933 3417 14967 3451
rect 19073 3349 19107 3383
rect 28641 2601 28675 2635
rect 1777 2397 1811 2431
rect 5457 2397 5491 2431
rect 17049 2397 17083 2431
rect 22753 2397 22787 2431
rect 30665 2397 30699 2431
rect 1409 2329 1443 2363
rect 10885 2329 10919 2363
rect 11253 2329 11287 2363
rect 28549 2329 28583 2363
rect 5365 2261 5399 2295
rect 16773 2261 16807 2295
rect 22845 2261 22879 2295
rect 30849 2261 30883 2295
<< metal1 >>
rect 1104 32122 31280 32144
rect 1104 32070 4182 32122
rect 4234 32070 4246 32122
rect 4298 32070 4310 32122
rect 4362 32070 4374 32122
rect 4426 32070 4438 32122
rect 4490 32070 4502 32122
rect 4554 32070 10182 32122
rect 10234 32070 10246 32122
rect 10298 32070 10310 32122
rect 10362 32070 10374 32122
rect 10426 32070 10438 32122
rect 10490 32070 10502 32122
rect 10554 32070 16182 32122
rect 16234 32070 16246 32122
rect 16298 32070 16310 32122
rect 16362 32070 16374 32122
rect 16426 32070 16438 32122
rect 16490 32070 16502 32122
rect 16554 32070 22182 32122
rect 22234 32070 22246 32122
rect 22298 32070 22310 32122
rect 22362 32070 22374 32122
rect 22426 32070 22438 32122
rect 22490 32070 22502 32122
rect 22554 32070 28182 32122
rect 28234 32070 28246 32122
rect 28298 32070 28310 32122
rect 28362 32070 28374 32122
rect 28426 32070 28438 32122
rect 28490 32070 28502 32122
rect 28554 32070 31280 32122
rect 1104 32048 31280 32070
rect 17865 32011 17923 32017
rect 17865 31977 17877 32011
rect 17911 32008 17923 32011
rect 18046 32008 18052 32020
rect 17911 31980 18052 32008
rect 17911 31977 17923 31980
rect 17865 31971 17923 31977
rect 18046 31968 18052 31980
rect 18104 31968 18110 32020
rect 23842 31968 23848 32020
rect 23900 32008 23906 32020
rect 24581 32011 24639 32017
rect 24581 32008 24593 32011
rect 23900 31980 24593 32008
rect 23900 31968 23906 31980
rect 24581 31977 24593 31980
rect 24627 31977 24639 32011
rect 24581 31971 24639 31977
rect 7561 31943 7619 31949
rect 7561 31909 7573 31943
rect 7607 31940 7619 31943
rect 18782 31940 18788 31952
rect 7607 31912 18788 31940
rect 7607 31909 7619 31912
rect 7561 31903 7619 31909
rect 18782 31900 18788 31912
rect 18840 31900 18846 31952
rect 1302 31764 1308 31816
rect 1360 31804 1366 31816
rect 1489 31807 1547 31813
rect 1489 31804 1501 31807
rect 1360 31776 1501 31804
rect 1360 31764 1366 31776
rect 1489 31773 1501 31776
rect 1535 31773 1547 31807
rect 1489 31767 1547 31773
rect 1670 31764 1676 31816
rect 1728 31764 1734 31816
rect 7098 31764 7104 31816
rect 7156 31804 7162 31816
rect 7285 31807 7343 31813
rect 7285 31804 7297 31807
rect 7156 31776 7297 31804
rect 7156 31764 7162 31776
rect 7285 31773 7297 31776
rect 7331 31773 7343 31807
rect 7285 31767 7343 31773
rect 12250 31764 12256 31816
rect 12308 31804 12314 31816
rect 12345 31807 12403 31813
rect 12345 31804 12357 31807
rect 12308 31776 12357 31804
rect 12308 31764 12314 31776
rect 12345 31773 12357 31776
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 18138 31764 18144 31816
rect 18196 31764 18202 31816
rect 18874 31764 18880 31816
rect 18932 31764 18938 31816
rect 24486 31764 24492 31816
rect 24544 31764 24550 31816
rect 29638 31764 29644 31816
rect 29696 31804 29702 31816
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29696 31776 29745 31804
rect 29696 31764 29702 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29733 31767 29791 31773
rect 12526 31628 12532 31680
rect 12584 31628 12590 31680
rect 18322 31628 18328 31680
rect 18380 31628 18386 31680
rect 26694 31628 26700 31680
rect 26752 31668 26758 31680
rect 29917 31671 29975 31677
rect 29917 31668 29929 31671
rect 26752 31640 29929 31668
rect 26752 31628 26758 31640
rect 29917 31637 29929 31640
rect 29963 31637 29975 31671
rect 29917 31631 29975 31637
rect 1104 31578 31280 31600
rect 1104 31526 4922 31578
rect 4974 31526 4986 31578
rect 5038 31526 5050 31578
rect 5102 31526 5114 31578
rect 5166 31526 5178 31578
rect 5230 31526 5242 31578
rect 5294 31526 10922 31578
rect 10974 31526 10986 31578
rect 11038 31526 11050 31578
rect 11102 31526 11114 31578
rect 11166 31526 11178 31578
rect 11230 31526 11242 31578
rect 11294 31526 16922 31578
rect 16974 31526 16986 31578
rect 17038 31526 17050 31578
rect 17102 31526 17114 31578
rect 17166 31526 17178 31578
rect 17230 31526 17242 31578
rect 17294 31526 22922 31578
rect 22974 31526 22986 31578
rect 23038 31526 23050 31578
rect 23102 31526 23114 31578
rect 23166 31526 23178 31578
rect 23230 31526 23242 31578
rect 23294 31526 28922 31578
rect 28974 31526 28986 31578
rect 29038 31526 29050 31578
rect 29102 31526 29114 31578
rect 29166 31526 29178 31578
rect 29230 31526 29242 31578
rect 29294 31526 31280 31578
rect 1104 31504 31280 31526
rect 11517 31467 11575 31473
rect 11517 31433 11529 31467
rect 11563 31433 11575 31467
rect 11517 31427 11575 31433
rect 17957 31467 18015 31473
rect 17957 31433 17969 31467
rect 18003 31464 18015 31467
rect 18322 31464 18328 31476
rect 18003 31436 18328 31464
rect 18003 31433 18015 31436
rect 17957 31427 18015 31433
rect 11149 31331 11207 31337
rect 11149 31297 11161 31331
rect 11195 31328 11207 31331
rect 11532 31328 11560 31427
rect 18322 31424 18328 31436
rect 18380 31424 18386 31476
rect 12526 31396 12532 31408
rect 11195 31300 11560 31328
rect 11808 31368 12532 31396
rect 11195 31297 11207 31300
rect 11149 31291 11207 31297
rect 7653 31263 7711 31269
rect 7653 31229 7665 31263
rect 7699 31260 7711 31263
rect 8570 31260 8576 31272
rect 7699 31232 8576 31260
rect 7699 31229 7711 31232
rect 7653 31223 7711 31229
rect 8570 31220 8576 31232
rect 8628 31220 8634 31272
rect 9122 31220 9128 31272
rect 9180 31260 9186 31272
rect 11808 31260 11836 31368
rect 12526 31356 12532 31368
rect 12584 31356 12590 31408
rect 18049 31399 18107 31405
rect 18049 31365 18061 31399
rect 18095 31396 18107 31399
rect 21082 31396 21088 31408
rect 18095 31368 21088 31396
rect 18095 31365 18107 31368
rect 18049 31359 18107 31365
rect 21082 31356 21088 31368
rect 21140 31356 21146 31408
rect 11885 31331 11943 31337
rect 11885 31297 11897 31331
rect 11931 31328 11943 31331
rect 12345 31331 12403 31337
rect 12345 31328 12357 31331
rect 11931 31300 12357 31328
rect 11931 31297 11943 31300
rect 11885 31291 11943 31297
rect 12345 31297 12357 31300
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 18785 31331 18843 31337
rect 18785 31297 18797 31331
rect 18831 31328 18843 31331
rect 19245 31331 19303 31337
rect 19245 31328 19257 31331
rect 18831 31300 19257 31328
rect 18831 31297 18843 31300
rect 18785 31291 18843 31297
rect 19245 31297 19257 31300
rect 19291 31297 19303 31331
rect 19245 31291 19303 31297
rect 20714 31288 20720 31340
rect 20772 31288 20778 31340
rect 21358 31288 21364 31340
rect 21416 31288 21422 31340
rect 23845 31331 23903 31337
rect 23845 31297 23857 31331
rect 23891 31328 23903 31331
rect 24210 31328 24216 31340
rect 23891 31300 24216 31328
rect 23891 31297 23903 31300
rect 23845 31291 23903 31297
rect 24210 31288 24216 31300
rect 24268 31288 24274 31340
rect 11977 31263 12035 31269
rect 11977 31260 11989 31263
rect 9180 31232 11989 31260
rect 9180 31220 9186 31232
rect 11977 31229 11989 31232
rect 12023 31229 12035 31263
rect 11977 31223 12035 31229
rect 12161 31263 12219 31269
rect 12161 31229 12173 31263
rect 12207 31229 12219 31263
rect 12161 31223 12219 31229
rect 12176 31192 12204 31223
rect 12894 31220 12900 31272
rect 12952 31220 12958 31272
rect 17954 31220 17960 31272
rect 18012 31260 18018 31272
rect 18141 31263 18199 31269
rect 18141 31260 18153 31263
rect 18012 31232 18153 31260
rect 18012 31220 18018 31232
rect 18141 31229 18153 31232
rect 18187 31260 18199 31263
rect 18187 31232 18644 31260
rect 18187 31229 18199 31232
rect 18141 31223 18199 31229
rect 14550 31192 14556 31204
rect 12176 31164 14556 31192
rect 14550 31152 14556 31164
rect 14608 31152 14614 31204
rect 16942 31152 16948 31204
rect 17000 31192 17006 31204
rect 18417 31195 18475 31201
rect 18417 31192 18429 31195
rect 17000 31164 18429 31192
rect 17000 31152 17006 31164
rect 18417 31161 18429 31164
rect 18463 31161 18475 31195
rect 18616 31192 18644 31232
rect 18690 31220 18696 31272
rect 18748 31260 18754 31272
rect 18877 31263 18935 31269
rect 18877 31260 18889 31263
rect 18748 31232 18889 31260
rect 18748 31220 18754 31232
rect 18877 31229 18889 31232
rect 18923 31229 18935 31263
rect 18877 31223 18935 31229
rect 18969 31263 19027 31269
rect 18969 31229 18981 31263
rect 19015 31229 19027 31263
rect 18969 31223 19027 31229
rect 18984 31192 19012 31223
rect 19794 31220 19800 31272
rect 19852 31220 19858 31272
rect 21634 31220 21640 31272
rect 21692 31260 21698 31272
rect 22373 31263 22431 31269
rect 22373 31260 22385 31263
rect 21692 31232 22385 31260
rect 21692 31220 21698 31232
rect 22373 31229 22385 31232
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 23290 31220 23296 31272
rect 23348 31220 23354 31272
rect 24670 31220 24676 31272
rect 24728 31220 24734 31272
rect 18616 31164 19012 31192
rect 18417 31155 18475 31161
rect 7006 31084 7012 31136
rect 7064 31084 7070 31136
rect 10962 31084 10968 31136
rect 11020 31084 11026 31136
rect 17586 31084 17592 31136
rect 17644 31084 17650 31136
rect 20530 31084 20536 31136
rect 20588 31084 20594 31136
rect 21542 31084 21548 31136
rect 21600 31084 21606 31136
rect 21818 31084 21824 31136
rect 21876 31084 21882 31136
rect 22738 31084 22744 31136
rect 22796 31084 22802 31136
rect 24026 31084 24032 31136
rect 24084 31084 24090 31136
rect 24118 31084 24124 31136
rect 24176 31084 24182 31136
rect 1104 31034 31280 31056
rect 1104 30982 4182 31034
rect 4234 30982 4246 31034
rect 4298 30982 4310 31034
rect 4362 30982 4374 31034
rect 4426 30982 4438 31034
rect 4490 30982 4502 31034
rect 4554 30982 10182 31034
rect 10234 30982 10246 31034
rect 10298 30982 10310 31034
rect 10362 30982 10374 31034
rect 10426 30982 10438 31034
rect 10490 30982 10502 31034
rect 10554 30982 16182 31034
rect 16234 30982 16246 31034
rect 16298 30982 16310 31034
rect 16362 30982 16374 31034
rect 16426 30982 16438 31034
rect 16490 30982 16502 31034
rect 16554 30982 22182 31034
rect 22234 30982 22246 31034
rect 22298 30982 22310 31034
rect 22362 30982 22374 31034
rect 22426 30982 22438 31034
rect 22490 30982 22502 31034
rect 22554 30982 28182 31034
rect 28234 30982 28246 31034
rect 28298 30982 28310 31034
rect 28362 30982 28374 31034
rect 28426 30982 28438 31034
rect 28490 30982 28502 31034
rect 28554 30982 31280 31034
rect 1104 30960 31280 30982
rect 12069 30923 12127 30929
rect 12069 30889 12081 30923
rect 12115 30920 12127 30923
rect 12894 30920 12900 30932
rect 12115 30892 12900 30920
rect 12115 30889 12127 30892
rect 12069 30883 12127 30889
rect 12894 30880 12900 30892
rect 12952 30880 12958 30932
rect 16942 30880 16948 30932
rect 17000 30880 17006 30932
rect 17586 30920 17592 30932
rect 17052 30892 17592 30920
rect 10410 30852 10416 30864
rect 9600 30824 10416 30852
rect 9600 30793 9628 30824
rect 10410 30812 10416 30824
rect 10468 30812 10474 30864
rect 9585 30787 9643 30793
rect 9585 30753 9597 30787
rect 9631 30753 9643 30787
rect 9585 30747 9643 30753
rect 9674 30744 9680 30796
rect 9732 30784 9738 30796
rect 10689 30787 10747 30793
rect 10689 30784 10701 30787
rect 9732 30756 10701 30784
rect 9732 30744 9738 30756
rect 10689 30753 10701 30756
rect 10735 30753 10747 30787
rect 10689 30747 10747 30753
rect 13541 30787 13599 30793
rect 13541 30753 13553 30787
rect 13587 30784 13599 30787
rect 13587 30756 14136 30784
rect 13587 30753 13599 30756
rect 13541 30747 13599 30753
rect 5445 30719 5503 30725
rect 5445 30685 5457 30719
rect 5491 30716 5503 30719
rect 5626 30716 5632 30728
rect 5491 30688 5632 30716
rect 5491 30685 5503 30688
rect 5445 30679 5503 30685
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30716 5779 30719
rect 7374 30716 7380 30728
rect 5767 30688 7380 30716
rect 5767 30685 5779 30688
rect 5721 30679 5779 30685
rect 7374 30676 7380 30688
rect 7432 30676 7438 30728
rect 10042 30716 10048 30728
rect 8772 30688 10048 30716
rect 5966 30651 6024 30657
rect 5966 30648 5978 30651
rect 5644 30620 5978 30648
rect 5644 30589 5672 30620
rect 5966 30617 5978 30620
rect 6012 30617 6024 30651
rect 5966 30611 6024 30617
rect 7644 30651 7702 30657
rect 7644 30617 7656 30651
rect 7690 30648 7702 30651
rect 8110 30648 8116 30660
rect 7690 30620 8116 30648
rect 7690 30617 7702 30620
rect 7644 30611 7702 30617
rect 8110 30608 8116 30620
rect 8168 30608 8174 30660
rect 5629 30583 5687 30589
rect 5629 30549 5641 30583
rect 5675 30549 5687 30583
rect 5629 30543 5687 30549
rect 7101 30583 7159 30589
rect 7101 30549 7113 30583
rect 7147 30580 7159 30583
rect 8570 30580 8576 30592
rect 7147 30552 8576 30580
rect 7147 30549 7159 30552
rect 7101 30543 7159 30549
rect 8570 30540 8576 30552
rect 8628 30540 8634 30592
rect 8772 30589 8800 30688
rect 10042 30676 10048 30688
rect 10100 30716 10106 30728
rect 10962 30725 10968 30728
rect 10321 30719 10379 30725
rect 10321 30716 10333 30719
rect 10100 30688 10333 30716
rect 10100 30676 10106 30688
rect 10321 30685 10333 30688
rect 10367 30685 10379 30719
rect 10956 30716 10968 30725
rect 10923 30688 10968 30716
rect 10321 30679 10379 30685
rect 10956 30679 10968 30688
rect 10962 30676 10968 30679
rect 11020 30676 11026 30728
rect 13725 30719 13783 30725
rect 13725 30685 13737 30719
rect 13771 30716 13783 30719
rect 13998 30716 14004 30728
rect 13771 30688 14004 30716
rect 13771 30685 13783 30688
rect 13725 30679 13783 30685
rect 13998 30676 14004 30688
rect 14056 30676 14062 30728
rect 14108 30725 14136 30756
rect 14093 30719 14151 30725
rect 14093 30685 14105 30719
rect 14139 30716 14151 30719
rect 14642 30716 14648 30728
rect 14139 30688 14648 30716
rect 14139 30685 14151 30688
rect 14093 30679 14151 30685
rect 14642 30676 14648 30688
rect 14700 30676 14706 30728
rect 16117 30719 16175 30725
rect 16117 30716 16129 30719
rect 15488 30688 16129 30716
rect 9309 30651 9367 30657
rect 9309 30617 9321 30651
rect 9355 30648 9367 30651
rect 9769 30651 9827 30657
rect 9769 30648 9781 30651
rect 9355 30620 9781 30648
rect 9355 30617 9367 30620
rect 9309 30611 9367 30617
rect 9769 30617 9781 30620
rect 9815 30617 9827 30651
rect 9769 30611 9827 30617
rect 11882 30608 11888 30660
rect 11940 30648 11946 30660
rect 11940 30620 12388 30648
rect 11940 30608 11946 30620
rect 12360 30592 12388 30620
rect 12802 30608 12808 30660
rect 12860 30648 12866 30660
rect 13274 30651 13332 30657
rect 13274 30648 13286 30651
rect 12860 30620 13286 30648
rect 12860 30608 12866 30620
rect 13274 30617 13286 30620
rect 13320 30617 13332 30651
rect 14338 30651 14396 30657
rect 14338 30648 14350 30651
rect 13274 30611 13332 30617
rect 13924 30620 14350 30648
rect 8757 30583 8815 30589
rect 8757 30549 8769 30583
rect 8803 30549 8815 30583
rect 8757 30543 8815 30549
rect 8938 30540 8944 30592
rect 8996 30540 9002 30592
rect 9122 30540 9128 30592
rect 9180 30580 9186 30592
rect 9401 30583 9459 30589
rect 9401 30580 9413 30583
rect 9180 30552 9413 30580
rect 9180 30540 9186 30552
rect 9401 30549 9413 30552
rect 9447 30549 9459 30583
rect 9401 30543 9459 30549
rect 12066 30540 12072 30592
rect 12124 30580 12130 30592
rect 12161 30583 12219 30589
rect 12161 30580 12173 30583
rect 12124 30552 12173 30580
rect 12124 30540 12130 30552
rect 12161 30549 12173 30552
rect 12207 30549 12219 30583
rect 12161 30543 12219 30549
rect 12342 30540 12348 30592
rect 12400 30540 12406 30592
rect 13924 30589 13952 30620
rect 14338 30617 14350 30620
rect 14384 30617 14396 30651
rect 14338 30611 14396 30617
rect 13909 30583 13967 30589
rect 13909 30549 13921 30583
rect 13955 30549 13967 30583
rect 13909 30543 13967 30549
rect 15010 30540 15016 30592
rect 15068 30580 15074 30592
rect 15488 30589 15516 30688
rect 16117 30685 16129 30688
rect 16163 30685 16175 30719
rect 16117 30679 16175 30685
rect 16761 30719 16819 30725
rect 16761 30685 16773 30719
rect 16807 30716 16819 30719
rect 16960 30716 16988 30880
rect 17052 30725 17080 30892
rect 17586 30880 17592 30892
rect 17644 30880 17650 30932
rect 18693 30923 18751 30929
rect 18693 30889 18705 30923
rect 18739 30920 18751 30923
rect 19794 30920 19800 30932
rect 18739 30892 19800 30920
rect 18739 30889 18751 30892
rect 18693 30883 18751 30889
rect 19794 30880 19800 30892
rect 19852 30880 19858 30932
rect 21542 30880 21548 30932
rect 21600 30880 21606 30932
rect 22830 30880 22836 30932
rect 22888 30920 22894 30932
rect 23109 30923 23167 30929
rect 23109 30920 23121 30923
rect 22888 30892 23121 30920
rect 22888 30880 22894 30892
rect 23109 30889 23121 30892
rect 23155 30920 23167 30923
rect 23290 30920 23296 30932
rect 23155 30892 23296 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 23290 30880 23296 30892
rect 23348 30880 23354 30932
rect 24118 30880 24124 30932
rect 24176 30880 24182 30932
rect 24210 30880 24216 30932
rect 24268 30880 24274 30932
rect 24397 30923 24455 30929
rect 24397 30889 24409 30923
rect 24443 30920 24455 30923
rect 24670 30920 24676 30932
rect 24443 30892 24676 30920
rect 24443 30889 24455 30892
rect 24397 30883 24455 30889
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 21560 30784 21588 30880
rect 23661 30787 23719 30793
rect 21560 30756 21864 30784
rect 16807 30688 16988 30716
rect 17037 30719 17095 30725
rect 16807 30685 16819 30688
rect 16761 30679 16819 30685
rect 17037 30685 17049 30719
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 17310 30676 17316 30728
rect 17368 30676 17374 30728
rect 19978 30676 19984 30728
rect 20036 30716 20042 30728
rect 20257 30719 20315 30725
rect 20257 30716 20269 30719
rect 20036 30688 20269 30716
rect 20036 30676 20042 30688
rect 20257 30685 20269 30688
rect 20303 30716 20315 30719
rect 21729 30719 21787 30725
rect 21729 30716 21741 30719
rect 20303 30688 21741 30716
rect 20303 30685 20315 30688
rect 20257 30679 20315 30685
rect 21729 30685 21741 30688
rect 21775 30685 21787 30719
rect 21836 30716 21864 30756
rect 23661 30753 23673 30787
rect 23707 30753 23719 30787
rect 23661 30747 23719 30753
rect 21985 30719 22043 30725
rect 21985 30716 21997 30719
rect 21836 30688 21997 30716
rect 21729 30679 21787 30685
rect 21985 30685 21997 30688
rect 22031 30685 22043 30719
rect 21985 30679 22043 30685
rect 23676 30660 23704 30747
rect 23845 30719 23903 30725
rect 23845 30685 23857 30719
rect 23891 30716 23903 30719
rect 24136 30716 24164 30880
rect 23891 30688 24164 30716
rect 23891 30685 23903 30688
rect 23845 30679 23903 30685
rect 24946 30676 24952 30728
rect 25004 30716 25010 30728
rect 25777 30719 25835 30725
rect 25777 30716 25789 30719
rect 25004 30688 25789 30716
rect 25004 30676 25010 30688
rect 25777 30685 25789 30688
rect 25823 30685 25835 30719
rect 25777 30679 25835 30685
rect 20530 30657 20536 30660
rect 17558 30651 17616 30657
rect 17558 30648 17570 30651
rect 16960 30620 17570 30648
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15068 30552 15485 30580
rect 15068 30540 15074 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 15473 30543 15531 30549
rect 15562 30540 15568 30592
rect 15620 30540 15626 30592
rect 16960 30589 16988 30620
rect 17558 30617 17570 30620
rect 17604 30617 17616 30651
rect 20524 30648 20536 30657
rect 20491 30620 20536 30648
rect 17558 30611 17616 30617
rect 20524 30611 20536 30620
rect 20530 30608 20536 30611
rect 20588 30608 20594 30660
rect 21082 30608 21088 30660
rect 21140 30648 21146 30660
rect 21140 30620 22094 30648
rect 21140 30608 21146 30620
rect 16945 30583 17003 30589
rect 16945 30549 16957 30583
rect 16991 30549 17003 30583
rect 16945 30543 17003 30549
rect 17221 30583 17279 30589
rect 17221 30549 17233 30583
rect 17267 30580 17279 30583
rect 17402 30580 17408 30592
rect 17267 30552 17408 30580
rect 17267 30549 17279 30552
rect 17221 30543 17279 30549
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 21634 30540 21640 30592
rect 21692 30540 21698 30592
rect 22066 30580 22094 30620
rect 23658 30608 23664 30660
rect 23716 30608 23722 30660
rect 24026 30608 24032 30660
rect 24084 30648 24090 30660
rect 25510 30651 25568 30657
rect 25510 30648 25522 30651
rect 24084 30620 25522 30648
rect 24084 30608 24090 30620
rect 25510 30617 25522 30620
rect 25556 30617 25568 30651
rect 25510 30611 25568 30617
rect 23753 30583 23811 30589
rect 23753 30580 23765 30583
rect 22066 30552 23765 30580
rect 23753 30549 23765 30552
rect 23799 30580 23811 30583
rect 26694 30580 26700 30592
rect 23799 30552 26700 30580
rect 23799 30549 23811 30552
rect 23753 30543 23811 30549
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 1104 30490 31280 30512
rect 1104 30438 4922 30490
rect 4974 30438 4986 30490
rect 5038 30438 5050 30490
rect 5102 30438 5114 30490
rect 5166 30438 5178 30490
rect 5230 30438 5242 30490
rect 5294 30438 10922 30490
rect 10974 30438 10986 30490
rect 11038 30438 11050 30490
rect 11102 30438 11114 30490
rect 11166 30438 11178 30490
rect 11230 30438 11242 30490
rect 11294 30438 16922 30490
rect 16974 30438 16986 30490
rect 17038 30438 17050 30490
rect 17102 30438 17114 30490
rect 17166 30438 17178 30490
rect 17230 30438 17242 30490
rect 17294 30438 22922 30490
rect 22974 30438 22986 30490
rect 23038 30438 23050 30490
rect 23102 30438 23114 30490
rect 23166 30438 23178 30490
rect 23230 30438 23242 30490
rect 23294 30438 28922 30490
rect 28974 30438 28986 30490
rect 29038 30438 29050 30490
rect 29102 30438 29114 30490
rect 29166 30438 29178 30490
rect 29230 30438 29242 30490
rect 29294 30438 31280 30490
rect 1104 30416 31280 30438
rect 5626 30336 5632 30388
rect 5684 30376 5690 30388
rect 6365 30379 6423 30385
rect 6365 30376 6377 30379
rect 5684 30348 6377 30376
rect 5684 30336 5690 30348
rect 6365 30345 6377 30348
rect 6411 30345 6423 30379
rect 6365 30339 6423 30345
rect 7006 30336 7012 30388
rect 7064 30336 7070 30388
rect 8110 30336 8116 30388
rect 8168 30336 8174 30388
rect 8938 30336 8944 30388
rect 8996 30336 9002 30388
rect 9646 30348 12020 30376
rect 6733 30311 6791 30317
rect 6733 30277 6745 30311
rect 6779 30308 6791 30311
rect 7024 30308 7052 30336
rect 6779 30280 7052 30308
rect 6779 30277 6791 30280
rect 6733 30271 6791 30277
rect 934 30200 940 30252
rect 992 30240 998 30252
rect 1397 30243 1455 30249
rect 1397 30240 1409 30243
rect 992 30212 1409 30240
rect 992 30200 998 30212
rect 1397 30209 1409 30212
rect 1443 30209 1455 30243
rect 8018 30240 8024 30252
rect 1397 30203 1455 30209
rect 6840 30212 8024 30240
rect 6840 30181 6868 30212
rect 8018 30200 8024 30212
rect 8076 30240 8082 30252
rect 8297 30243 8355 30249
rect 8076 30212 8248 30240
rect 8076 30200 8082 30212
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 1596 30144 6837 30172
rect 1596 30113 1624 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 6825 30135 6883 30141
rect 6917 30175 6975 30181
rect 6917 30141 6929 30175
rect 6963 30141 6975 30175
rect 8220 30172 8248 30212
rect 8297 30209 8309 30243
rect 8343 30240 8355 30243
rect 8956 30240 8984 30336
rect 9646 30308 9674 30348
rect 8343 30212 8984 30240
rect 9048 30280 9674 30308
rect 8343 30209 8355 30212
rect 8297 30203 8355 30209
rect 9048 30172 9076 30280
rect 11882 30268 11888 30320
rect 11940 30268 11946 30320
rect 11992 30317 12020 30348
rect 12250 30336 12256 30388
rect 12308 30376 12314 30388
rect 12308 30348 12434 30376
rect 12308 30336 12314 30348
rect 11977 30311 12035 30317
rect 11977 30277 11989 30311
rect 12023 30308 12035 30311
rect 12406 30308 12434 30348
rect 13998 30336 14004 30388
rect 14056 30336 14062 30388
rect 15562 30336 15568 30388
rect 15620 30336 15626 30388
rect 17402 30336 17408 30388
rect 17460 30336 17466 30388
rect 18690 30336 18696 30388
rect 18748 30376 18754 30388
rect 20625 30379 20683 30385
rect 18748 30348 19656 30376
rect 18748 30336 18754 30348
rect 14369 30311 14427 30317
rect 12023 30280 12204 30308
rect 12406 30280 12940 30308
rect 12023 30277 12035 30280
rect 11977 30271 12035 30277
rect 10965 30243 11023 30249
rect 10965 30209 10977 30243
rect 11011 30240 11023 30243
rect 11514 30240 11520 30252
rect 11011 30212 11520 30240
rect 11011 30209 11023 30212
rect 10965 30203 11023 30209
rect 11514 30200 11520 30212
rect 11572 30200 11578 30252
rect 8220 30144 9076 30172
rect 6917 30135 6975 30141
rect 1581 30107 1639 30113
rect 1581 30073 1593 30107
rect 1627 30073 1639 30107
rect 1581 30067 1639 30073
rect 5994 30064 6000 30116
rect 6052 30104 6058 30116
rect 6932 30104 6960 30135
rect 10410 30132 10416 30184
rect 10468 30172 10474 30184
rect 10778 30172 10784 30184
rect 10468 30144 10784 30172
rect 10468 30132 10474 30144
rect 10778 30132 10784 30144
rect 10836 30172 10842 30184
rect 12069 30175 12127 30181
rect 12069 30172 12081 30175
rect 10836 30144 12081 30172
rect 10836 30132 10842 30144
rect 12069 30141 12081 30144
rect 12115 30141 12127 30175
rect 12176 30172 12204 30280
rect 12342 30200 12348 30252
rect 12400 30200 12406 30252
rect 12912 30249 12940 30280
rect 14369 30277 14381 30311
rect 14415 30308 14427 30311
rect 15580 30308 15608 30336
rect 14415 30280 15608 30308
rect 14415 30277 14427 30280
rect 14369 30271 14427 30277
rect 12897 30243 12955 30249
rect 12897 30209 12909 30243
rect 12943 30209 12955 30243
rect 12897 30203 12955 30209
rect 17221 30243 17279 30249
rect 17221 30209 17233 30243
rect 17267 30240 17279 30243
rect 17310 30240 17316 30252
rect 17267 30212 17316 30240
rect 17267 30209 17279 30212
rect 17221 30203 17279 30209
rect 17310 30200 17316 30212
rect 17368 30200 17374 30252
rect 17420 30240 17448 30336
rect 17477 30243 17535 30249
rect 17477 30240 17489 30243
rect 17420 30212 17489 30240
rect 17477 30209 17489 30212
rect 17523 30209 17535 30243
rect 17477 30203 17535 30209
rect 14461 30175 14519 30181
rect 14461 30172 14473 30175
rect 12176 30144 14473 30172
rect 12069 30135 12127 30141
rect 14461 30141 14473 30144
rect 14507 30141 14519 30175
rect 14461 30135 14519 30141
rect 14550 30132 14556 30184
rect 14608 30132 14614 30184
rect 19628 30172 19656 30348
rect 20625 30345 20637 30379
rect 20671 30376 20683 30379
rect 20714 30376 20720 30388
rect 20671 30348 20720 30376
rect 20671 30345 20683 30348
rect 20625 30339 20683 30345
rect 20714 30336 20720 30348
rect 20772 30336 20778 30388
rect 20993 30379 21051 30385
rect 20993 30345 21005 30379
rect 21039 30376 21051 30379
rect 21818 30376 21824 30388
rect 21039 30348 21824 30376
rect 21039 30345 21051 30348
rect 20993 30339 21051 30345
rect 21818 30336 21824 30348
rect 21876 30336 21882 30388
rect 22189 30379 22247 30385
rect 22189 30345 22201 30379
rect 22235 30376 22247 30379
rect 22738 30376 22744 30388
rect 22235 30348 22744 30376
rect 22235 30345 22247 30348
rect 22189 30339 22247 30345
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 23124 30348 23336 30376
rect 19978 30268 19984 30320
rect 20036 30308 20042 30320
rect 23124 30308 23152 30348
rect 20036 30280 23152 30308
rect 23308 30308 23336 30348
rect 24946 30308 24952 30320
rect 23308 30280 24952 30308
rect 20036 30268 20042 30280
rect 21082 30200 21088 30252
rect 21140 30200 21146 30252
rect 22094 30240 22100 30252
rect 21192 30212 22100 30240
rect 21192 30172 21220 30212
rect 22094 30200 22100 30212
rect 22152 30240 22158 30252
rect 22281 30243 22339 30249
rect 22281 30240 22293 30243
rect 22152 30212 22293 30240
rect 22152 30200 22158 30212
rect 22281 30209 22293 30212
rect 22327 30209 22339 30243
rect 22281 30203 22339 30209
rect 23014 30200 23020 30252
rect 23072 30200 23078 30252
rect 23198 30240 23204 30252
rect 23124 30212 23204 30240
rect 19628 30144 21220 30172
rect 21269 30175 21327 30181
rect 21269 30141 21281 30175
rect 21315 30141 21327 30175
rect 21269 30135 21327 30141
rect 22465 30175 22523 30181
rect 22465 30141 22477 30175
rect 22511 30172 22523 30175
rect 23124 30172 23152 30212
rect 23198 30200 23204 30212
rect 23256 30200 23262 30252
rect 23308 30249 23336 30280
rect 24946 30268 24952 30280
rect 25004 30268 25010 30320
rect 23293 30243 23351 30249
rect 23293 30209 23305 30243
rect 23339 30209 23351 30243
rect 23549 30243 23607 30249
rect 23549 30240 23561 30243
rect 23293 30203 23351 30209
rect 23400 30212 23561 30240
rect 23400 30172 23428 30212
rect 23549 30209 23561 30212
rect 23595 30209 23607 30243
rect 23549 30203 23607 30209
rect 25317 30175 25375 30181
rect 25317 30172 25329 30175
rect 22511 30144 23152 30172
rect 23216 30144 23428 30172
rect 24688 30144 25329 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 6052 30076 6960 30104
rect 6052 30064 6058 30076
rect 11514 30064 11520 30116
rect 11572 30064 11578 30116
rect 12176 30076 12434 30104
rect 11149 30039 11207 30045
rect 11149 30005 11161 30039
rect 11195 30036 11207 30039
rect 12176 30036 12204 30076
rect 11195 30008 12204 30036
rect 12406 30036 12434 30076
rect 12802 30036 12808 30048
rect 12406 30008 12808 30036
rect 11195 30005 11207 30008
rect 11149 29999 11207 30005
rect 12802 29996 12808 30008
rect 12860 29996 12866 30048
rect 14568 30036 14596 30132
rect 18601 30107 18659 30113
rect 18601 30073 18613 30107
rect 18647 30104 18659 30107
rect 18874 30104 18880 30116
rect 18647 30076 18880 30104
rect 18647 30073 18659 30076
rect 18601 30067 18659 30073
rect 18874 30064 18880 30076
rect 18932 30064 18938 30116
rect 17954 30036 17960 30048
rect 14568 30008 17960 30036
rect 17954 29996 17960 30008
rect 18012 29996 18018 30048
rect 20898 29996 20904 30048
rect 20956 30036 20962 30048
rect 21284 30036 21312 30135
rect 23216 30113 23244 30144
rect 23201 30107 23259 30113
rect 23201 30073 23213 30107
rect 23247 30073 23259 30107
rect 23201 30067 23259 30073
rect 20956 30008 21312 30036
rect 20956 29996 20962 30008
rect 21358 29996 21364 30048
rect 21416 30036 21422 30048
rect 21821 30039 21879 30045
rect 21821 30036 21833 30039
rect 21416 30008 21833 30036
rect 21416 29996 21422 30008
rect 21821 30005 21833 30008
rect 21867 30005 21879 30039
rect 21821 29999 21879 30005
rect 23106 29996 23112 30048
rect 23164 30036 23170 30048
rect 24688 30045 24716 30144
rect 25317 30141 25329 30144
rect 25363 30141 25375 30175
rect 25317 30135 25375 30141
rect 24673 30039 24731 30045
rect 24673 30036 24685 30039
rect 23164 30008 24685 30036
rect 23164 29996 23170 30008
rect 24673 30005 24685 30008
rect 24719 30005 24731 30039
rect 24673 29999 24731 30005
rect 24762 29996 24768 30048
rect 24820 29996 24826 30048
rect 1104 29946 31280 29968
rect 1104 29894 4182 29946
rect 4234 29894 4246 29946
rect 4298 29894 4310 29946
rect 4362 29894 4374 29946
rect 4426 29894 4438 29946
rect 4490 29894 4502 29946
rect 4554 29894 10182 29946
rect 10234 29894 10246 29946
rect 10298 29894 10310 29946
rect 10362 29894 10374 29946
rect 10426 29894 10438 29946
rect 10490 29894 10502 29946
rect 10554 29894 16182 29946
rect 16234 29894 16246 29946
rect 16298 29894 16310 29946
rect 16362 29894 16374 29946
rect 16426 29894 16438 29946
rect 16490 29894 16502 29946
rect 16554 29894 22182 29946
rect 22234 29894 22246 29946
rect 22298 29894 22310 29946
rect 22362 29894 22374 29946
rect 22426 29894 22438 29946
rect 22490 29894 22502 29946
rect 22554 29894 28182 29946
rect 28234 29894 28246 29946
rect 28298 29894 28310 29946
rect 28362 29894 28374 29946
rect 28426 29894 28438 29946
rect 28490 29894 28502 29946
rect 28554 29894 31280 29946
rect 1104 29872 31280 29894
rect 11974 29792 11980 29844
rect 12032 29832 12038 29844
rect 15286 29832 15292 29844
rect 12032 29804 15292 29832
rect 12032 29792 12038 29804
rect 15286 29792 15292 29804
rect 15344 29792 15350 29844
rect 23014 29792 23020 29844
rect 23072 29832 23078 29844
rect 23477 29835 23535 29841
rect 23477 29832 23489 29835
rect 23072 29804 23489 29832
rect 23072 29792 23078 29804
rect 23477 29801 23489 29804
rect 23523 29801 23535 29835
rect 23477 29795 23535 29801
rect 24762 29792 24768 29844
rect 24820 29792 24826 29844
rect 19981 29767 20039 29773
rect 19981 29733 19993 29767
rect 20027 29764 20039 29767
rect 21910 29764 21916 29776
rect 20027 29736 21916 29764
rect 20027 29733 20039 29736
rect 19981 29727 20039 29733
rect 21910 29724 21916 29736
rect 21968 29724 21974 29776
rect 23934 29764 23940 29776
rect 23032 29736 23940 29764
rect 9968 29668 10456 29696
rect 8478 29588 8484 29640
rect 8536 29588 8542 29640
rect 9968 29637 9996 29668
rect 9953 29631 10011 29637
rect 9953 29628 9965 29631
rect 9324 29600 9965 29628
rect 9324 29504 9352 29600
rect 9953 29597 9965 29600
rect 9999 29597 10011 29631
rect 9953 29591 10011 29597
rect 10042 29588 10048 29640
rect 10100 29628 10106 29640
rect 10428 29637 10456 29668
rect 10137 29631 10195 29637
rect 10137 29628 10149 29631
rect 10100 29600 10149 29628
rect 10100 29588 10106 29600
rect 10137 29597 10149 29600
rect 10183 29597 10195 29631
rect 10137 29591 10195 29597
rect 10413 29631 10471 29637
rect 10413 29597 10425 29631
rect 10459 29597 10471 29631
rect 10413 29591 10471 29597
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 11330 29628 11336 29640
rect 10551 29600 11336 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 11330 29588 11336 29600
rect 11388 29588 11394 29640
rect 12342 29588 12348 29640
rect 12400 29588 12406 29640
rect 14642 29588 14648 29640
rect 14700 29628 14706 29640
rect 14700 29600 15884 29628
rect 14700 29588 14706 29600
rect 10321 29563 10379 29569
rect 10321 29529 10333 29563
rect 10367 29560 10379 29563
rect 12250 29560 12256 29572
rect 10367 29532 12256 29560
rect 10367 29529 10379 29532
rect 10321 29523 10379 29529
rect 12250 29520 12256 29532
rect 12308 29520 12314 29572
rect 14918 29569 14924 29572
rect 14912 29523 14924 29569
rect 14918 29520 14924 29523
rect 14976 29520 14982 29572
rect 15378 29560 15384 29572
rect 15028 29532 15384 29560
rect 8294 29452 8300 29504
rect 8352 29452 8358 29504
rect 9306 29452 9312 29504
rect 9364 29452 9370 29504
rect 9398 29452 9404 29504
rect 9456 29452 9462 29504
rect 10686 29452 10692 29504
rect 10744 29452 10750 29504
rect 11698 29452 11704 29504
rect 11756 29452 11762 29504
rect 12526 29452 12532 29504
rect 12584 29492 12590 29504
rect 15028 29492 15056 29532
rect 15378 29520 15384 29532
rect 15436 29520 15442 29572
rect 15856 29560 15884 29600
rect 16022 29588 16028 29640
rect 16080 29628 16086 29640
rect 16669 29631 16727 29637
rect 16669 29628 16681 29631
rect 16080 29600 16681 29628
rect 16080 29588 16086 29600
rect 16669 29597 16681 29600
rect 16715 29597 16727 29631
rect 16669 29591 16727 29597
rect 17310 29588 17316 29640
rect 17368 29588 17374 29640
rect 18874 29588 18880 29640
rect 18932 29628 18938 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 18932 29600 19441 29628
rect 18932 29588 18938 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19705 29631 19763 29637
rect 19705 29628 19717 29631
rect 19429 29591 19487 29597
rect 19536 29600 19717 29628
rect 17328 29560 17356 29588
rect 15856 29532 17356 29560
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 19536 29560 19564 29600
rect 19705 29597 19717 29600
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29628 19855 29631
rect 19886 29628 19892 29640
rect 19843 29600 19892 29628
rect 19843 29597 19855 29600
rect 19797 29591 19855 29597
rect 19886 29588 19892 29600
rect 19944 29588 19950 29640
rect 20990 29588 20996 29640
rect 21048 29588 21054 29640
rect 22830 29588 22836 29640
rect 22888 29588 22894 29640
rect 23032 29637 23060 29736
rect 23934 29724 23940 29736
rect 23992 29764 23998 29776
rect 24394 29764 24400 29776
rect 23992 29736 24400 29764
rect 23992 29724 23998 29736
rect 24394 29724 24400 29736
rect 24452 29724 24458 29776
rect 24121 29699 24179 29705
rect 24121 29665 24133 29699
rect 24167 29696 24179 29699
rect 24486 29696 24492 29708
rect 24167 29668 24492 29696
rect 24167 29665 24179 29668
rect 24121 29659 24179 29665
rect 24486 29656 24492 29668
rect 24544 29656 24550 29708
rect 23017 29631 23075 29637
rect 23017 29597 23029 29631
rect 23063 29597 23075 29631
rect 23017 29591 23075 29597
rect 23106 29588 23112 29640
rect 23164 29588 23170 29640
rect 23201 29631 23259 29637
rect 23201 29597 23213 29631
rect 23247 29597 23259 29631
rect 23201 29591 23259 29597
rect 23845 29631 23903 29637
rect 23845 29597 23857 29631
rect 23891 29628 23903 29631
rect 24780 29628 24808 29792
rect 24946 29656 24952 29708
rect 25004 29656 25010 29708
rect 23891 29600 24808 29628
rect 24964 29628 24992 29656
rect 25961 29631 26019 29637
rect 25961 29628 25973 29631
rect 24964 29600 25973 29628
rect 23891 29597 23903 29600
rect 23845 29591 23903 29597
rect 25961 29597 25973 29600
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 19392 29532 19564 29560
rect 19392 29520 19398 29532
rect 19610 29520 19616 29572
rect 19668 29520 19674 29572
rect 23216 29560 23244 29591
rect 25716 29563 25774 29569
rect 23216 29532 24348 29560
rect 24320 29504 24348 29532
rect 25716 29529 25728 29563
rect 25762 29560 25774 29563
rect 26234 29560 26240 29572
rect 25762 29532 26240 29560
rect 25762 29529 25774 29532
rect 25716 29523 25774 29529
rect 26234 29520 26240 29532
rect 26292 29520 26298 29572
rect 12584 29464 15056 29492
rect 12584 29452 12590 29464
rect 15194 29452 15200 29504
rect 15252 29492 15258 29504
rect 16022 29492 16028 29504
rect 15252 29464 16028 29492
rect 15252 29452 15258 29464
rect 16022 29452 16028 29464
rect 16080 29452 16086 29504
rect 16114 29452 16120 29504
rect 16172 29452 16178 29504
rect 20806 29452 20812 29504
rect 20864 29452 20870 29504
rect 23382 29452 23388 29504
rect 23440 29452 23446 29504
rect 23842 29452 23848 29504
rect 23900 29492 23906 29504
rect 23937 29495 23995 29501
rect 23937 29492 23949 29495
rect 23900 29464 23949 29492
rect 23900 29452 23906 29464
rect 23937 29461 23949 29464
rect 23983 29461 23995 29495
rect 23937 29455 23995 29461
rect 24302 29452 24308 29504
rect 24360 29452 24366 29504
rect 24578 29452 24584 29504
rect 24636 29452 24642 29504
rect 1104 29402 31280 29424
rect 1104 29350 4922 29402
rect 4974 29350 4986 29402
rect 5038 29350 5050 29402
rect 5102 29350 5114 29402
rect 5166 29350 5178 29402
rect 5230 29350 5242 29402
rect 5294 29350 10922 29402
rect 10974 29350 10986 29402
rect 11038 29350 11050 29402
rect 11102 29350 11114 29402
rect 11166 29350 11178 29402
rect 11230 29350 11242 29402
rect 11294 29350 16922 29402
rect 16974 29350 16986 29402
rect 17038 29350 17050 29402
rect 17102 29350 17114 29402
rect 17166 29350 17178 29402
rect 17230 29350 17242 29402
rect 17294 29350 22922 29402
rect 22974 29350 22986 29402
rect 23038 29350 23050 29402
rect 23102 29350 23114 29402
rect 23166 29350 23178 29402
rect 23230 29350 23242 29402
rect 23294 29350 28922 29402
rect 28974 29350 28986 29402
rect 29038 29350 29050 29402
rect 29102 29350 29114 29402
rect 29166 29350 29178 29402
rect 29230 29350 29242 29402
rect 29294 29350 31280 29402
rect 1104 29328 31280 29350
rect 8294 29248 8300 29300
rect 8352 29248 8358 29300
rect 9306 29248 9312 29300
rect 9364 29248 9370 29300
rect 11698 29248 11704 29300
rect 11756 29288 11762 29300
rect 11885 29291 11943 29297
rect 11885 29288 11897 29291
rect 11756 29260 11897 29288
rect 11756 29248 11762 29260
rect 11885 29257 11897 29260
rect 11931 29257 11943 29291
rect 11885 29251 11943 29257
rect 12526 29248 12532 29300
rect 12584 29248 12590 29300
rect 14458 29288 14464 29300
rect 12636 29260 14464 29288
rect 8196 29223 8254 29229
rect 8196 29189 8208 29223
rect 8242 29220 8254 29223
rect 8312 29220 8340 29248
rect 8242 29192 8340 29220
rect 8242 29189 8254 29192
rect 8196 29183 8254 29189
rect 6549 29155 6607 29161
rect 6549 29121 6561 29155
rect 6595 29152 6607 29155
rect 7006 29152 7012 29164
rect 6595 29124 7012 29152
rect 6595 29121 6607 29124
rect 6549 29115 6607 29121
rect 7006 29112 7012 29124
rect 7064 29112 7070 29164
rect 7374 29112 7380 29164
rect 7432 29152 7438 29164
rect 7929 29155 7987 29161
rect 7929 29152 7941 29155
rect 7432 29124 7941 29152
rect 7432 29112 7438 29124
rect 7929 29121 7941 29124
rect 7975 29121 7987 29155
rect 7929 29115 7987 29121
rect 10220 29155 10278 29161
rect 10220 29121 10232 29155
rect 10266 29152 10278 29155
rect 10594 29152 10600 29164
rect 10266 29124 10600 29152
rect 10266 29121 10278 29124
rect 10220 29115 10278 29121
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 12544 29161 12572 29248
rect 12636 29229 12664 29260
rect 14458 29248 14464 29260
rect 14516 29248 14522 29300
rect 14642 29248 14648 29300
rect 14700 29248 14706 29300
rect 14829 29291 14887 29297
rect 14829 29257 14841 29291
rect 14875 29288 14887 29291
rect 14918 29288 14924 29300
rect 14875 29260 14924 29288
rect 14875 29257 14887 29260
rect 14829 29251 14887 29257
rect 14918 29248 14924 29260
rect 14976 29248 14982 29300
rect 15013 29291 15071 29297
rect 15013 29257 15025 29291
rect 15059 29257 15071 29291
rect 15013 29251 15071 29257
rect 12621 29223 12679 29229
rect 12621 29189 12633 29223
rect 12667 29189 12679 29223
rect 14660 29220 14688 29248
rect 12621 29183 12679 29189
rect 13096 29192 14688 29220
rect 12529 29155 12587 29161
rect 12529 29121 12541 29155
rect 12575 29121 12587 29155
rect 12529 29115 12587 29121
rect 12713 29155 12771 29161
rect 12713 29121 12725 29155
rect 12759 29121 12771 29155
rect 12713 29115 12771 29121
rect 6086 29044 6092 29096
rect 6144 29044 6150 29096
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 9953 29087 10011 29093
rect 9953 29084 9965 29087
rect 9732 29056 9965 29084
rect 9732 29044 9738 29056
rect 9953 29053 9965 29056
rect 9999 29053 10011 29087
rect 9953 29047 10011 29053
rect 11974 29044 11980 29096
rect 12032 29044 12038 29096
rect 12158 29044 12164 29096
rect 12216 29044 12222 29096
rect 12342 29044 12348 29096
rect 12400 29044 12406 29096
rect 11333 29019 11391 29025
rect 11333 28985 11345 29019
rect 11379 29016 11391 29019
rect 12360 29016 12388 29044
rect 11379 28988 12388 29016
rect 12728 29016 12756 29115
rect 12894 29112 12900 29164
rect 12952 29112 12958 29164
rect 13096 29161 13124 29192
rect 13081 29155 13139 29161
rect 13081 29121 13093 29155
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13170 29112 13176 29164
rect 13228 29152 13234 29164
rect 13337 29155 13395 29161
rect 13337 29152 13349 29155
rect 13228 29124 13349 29152
rect 13228 29112 13234 29124
rect 13337 29121 13349 29124
rect 13383 29121 13395 29155
rect 13337 29115 13395 29121
rect 14645 29155 14703 29161
rect 14645 29121 14657 29155
rect 14691 29152 14703 29155
rect 15028 29152 15056 29251
rect 15286 29248 15292 29300
rect 15344 29248 15350 29300
rect 15381 29291 15439 29297
rect 15381 29257 15393 29291
rect 15427 29288 15439 29291
rect 16114 29288 16120 29300
rect 15427 29260 16120 29288
rect 15427 29257 15439 29260
rect 15381 29251 15439 29257
rect 16114 29248 16120 29260
rect 16172 29248 16178 29300
rect 17957 29291 18015 29297
rect 17957 29257 17969 29291
rect 18003 29257 18015 29291
rect 19794 29288 19800 29300
rect 17957 29251 18015 29257
rect 19536 29260 19800 29288
rect 15304 29220 15332 29248
rect 15473 29223 15531 29229
rect 15473 29220 15485 29223
rect 15304 29192 15485 29220
rect 15473 29189 15485 29192
rect 15519 29189 15531 29223
rect 15473 29183 15531 29189
rect 14691 29124 15056 29152
rect 17865 29155 17923 29161
rect 14691 29121 14703 29124
rect 14645 29115 14703 29121
rect 17865 29121 17877 29155
rect 17911 29152 17923 29155
rect 17972 29152 18000 29251
rect 18417 29223 18475 29229
rect 18417 29189 18429 29223
rect 18463 29220 18475 29223
rect 19426 29220 19432 29232
rect 18463 29192 19432 29220
rect 18463 29189 18475 29192
rect 18417 29183 18475 29189
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 19536 29161 19564 29260
rect 19794 29248 19800 29260
rect 19852 29248 19858 29300
rect 20073 29291 20131 29297
rect 20073 29257 20085 29291
rect 20119 29288 20131 29291
rect 20714 29288 20720 29300
rect 20119 29260 20720 29288
rect 20119 29257 20131 29260
rect 20073 29251 20131 29257
rect 20714 29248 20720 29260
rect 20772 29248 20778 29300
rect 20806 29248 20812 29300
rect 20864 29248 20870 29300
rect 24578 29248 24584 29300
rect 24636 29248 24642 29300
rect 26234 29248 26240 29300
rect 26292 29248 26298 29300
rect 19610 29180 19616 29232
rect 19668 29220 19674 29232
rect 19705 29223 19763 29229
rect 19705 29220 19717 29223
rect 19668 29192 19717 29220
rect 19668 29180 19674 29192
rect 19705 29189 19717 29192
rect 19751 29189 19763 29223
rect 19705 29183 19763 29189
rect 20524 29223 20582 29229
rect 20524 29189 20536 29223
rect 20570 29220 20582 29223
rect 20824 29220 20852 29248
rect 20570 29192 20852 29220
rect 24305 29223 24363 29229
rect 20570 29189 20582 29192
rect 20524 29183 20582 29189
rect 24305 29189 24317 29223
rect 24351 29220 24363 29223
rect 24596 29220 24624 29248
rect 24351 29192 26096 29220
rect 24351 29189 24363 29192
rect 24305 29183 24363 29189
rect 17911 29124 18000 29152
rect 18325 29155 18383 29161
rect 17911 29121 17923 29124
rect 17865 29115 17923 29121
rect 18325 29121 18337 29155
rect 18371 29152 18383 29155
rect 18785 29155 18843 29161
rect 18785 29152 18797 29155
rect 18371 29124 18797 29152
rect 18371 29121 18383 29124
rect 18325 29115 18383 29121
rect 18785 29121 18797 29124
rect 18831 29121 18843 29155
rect 18785 29115 18843 29121
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 19794 29112 19800 29164
rect 19852 29112 19858 29164
rect 19886 29112 19892 29164
rect 19944 29152 19950 29164
rect 20346 29152 20352 29164
rect 19944 29124 20352 29152
rect 19944 29112 19950 29124
rect 20346 29112 20352 29124
rect 20404 29112 20410 29164
rect 24213 29155 24271 29161
rect 24213 29121 24225 29155
rect 24259 29152 24271 29155
rect 24259 29124 24348 29152
rect 24259 29121 24271 29124
rect 24213 29115 24271 29121
rect 15657 29087 15715 29093
rect 15657 29053 15669 29087
rect 15703 29084 15715 29087
rect 18601 29087 18659 29093
rect 18601 29084 18613 29087
rect 15703 29056 18613 29084
rect 15703 29053 15715 29056
rect 15657 29047 15715 29053
rect 18601 29053 18613 29056
rect 18647 29084 18659 29087
rect 18874 29084 18880 29096
rect 18647 29056 18880 29084
rect 18647 29053 18659 29056
rect 18601 29047 18659 29053
rect 18874 29044 18880 29056
rect 18932 29044 18938 29096
rect 19334 29044 19340 29096
rect 19392 29044 19398 29096
rect 19978 29044 19984 29096
rect 20036 29084 20042 29096
rect 20257 29087 20315 29093
rect 20257 29084 20269 29087
rect 20036 29056 20269 29084
rect 20036 29044 20042 29056
rect 20257 29053 20269 29056
rect 20303 29053 20315 29087
rect 22465 29087 22523 29093
rect 22465 29084 22477 29087
rect 20257 29047 20315 29053
rect 22066 29056 22477 29084
rect 21637 29019 21695 29025
rect 12728 28988 13124 29016
rect 11379 28985 11391 28988
rect 11333 28979 11391 28985
rect 13096 28960 13124 28988
rect 21637 28985 21649 29019
rect 21683 29016 21695 29019
rect 22066 29016 22094 29056
rect 22465 29053 22477 29056
rect 22511 29084 22523 29087
rect 22830 29084 22836 29096
rect 22511 29056 22836 29084
rect 22511 29053 22523 29056
rect 22465 29047 22523 29053
rect 22830 29044 22836 29056
rect 22888 29044 22894 29096
rect 24320 29028 24348 29124
rect 24394 29112 24400 29164
rect 24452 29112 24458 29164
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29152 24639 29155
rect 24670 29152 24676 29164
rect 24627 29124 24676 29152
rect 24627 29121 24639 29124
rect 24581 29115 24639 29121
rect 24670 29112 24676 29124
rect 24728 29112 24734 29164
rect 26068 29161 26096 29192
rect 25041 29155 25099 29161
rect 25041 29121 25053 29155
rect 25087 29152 25099 29155
rect 25501 29155 25559 29161
rect 25501 29152 25513 29155
rect 25087 29124 25513 29152
rect 25087 29121 25099 29124
rect 25041 29115 25099 29121
rect 25501 29121 25513 29124
rect 25547 29121 25559 29155
rect 25501 29115 25559 29121
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29121 26111 29155
rect 26053 29115 26111 29121
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 24486 29044 24492 29096
rect 24544 29084 24550 29096
rect 24765 29087 24823 29093
rect 24765 29084 24777 29087
rect 24544 29056 24777 29084
rect 24544 29044 24550 29056
rect 24688 29028 24716 29056
rect 24765 29053 24777 29056
rect 24811 29053 24823 29087
rect 24765 29047 24823 29053
rect 24946 29044 24952 29096
rect 25004 29044 25010 29096
rect 21683 28988 22094 29016
rect 21683 28985 21695 28988
rect 21637 28979 21695 28985
rect 24302 28976 24308 29028
rect 24360 28976 24366 29028
rect 24670 28976 24676 29028
rect 24728 28976 24734 29028
rect 25409 29019 25467 29025
rect 25409 28985 25421 29019
rect 25455 29016 25467 29019
rect 26436 29016 26464 29115
rect 25455 28988 26464 29016
rect 25455 28985 25467 28988
rect 25409 28979 25467 28985
rect 5534 28908 5540 28960
rect 5592 28908 5598 28960
rect 6362 28908 6368 28960
rect 6420 28908 6426 28960
rect 6454 28908 6460 28960
rect 6512 28948 6518 28960
rect 9122 28948 9128 28960
rect 6512 28920 9128 28948
rect 6512 28908 6518 28920
rect 9122 28908 9128 28920
rect 9180 28908 9186 28960
rect 11514 28908 11520 28960
rect 11572 28908 11578 28960
rect 11606 28908 11612 28960
rect 11664 28948 11670 28960
rect 12345 28951 12403 28957
rect 12345 28948 12357 28951
rect 11664 28920 12357 28948
rect 11664 28908 11670 28920
rect 12345 28917 12357 28920
rect 12391 28917 12403 28951
rect 12345 28911 12403 28917
rect 13078 28908 13084 28960
rect 13136 28948 13142 28960
rect 15102 28948 15108 28960
rect 13136 28920 15108 28948
rect 13136 28908 13142 28920
rect 15102 28908 15108 28920
rect 15160 28908 15166 28960
rect 17678 28908 17684 28960
rect 17736 28908 17742 28960
rect 21818 28908 21824 28960
rect 21876 28908 21882 28960
rect 24026 28908 24032 28960
rect 24084 28908 24090 28960
rect 1104 28858 31280 28880
rect 1104 28806 4182 28858
rect 4234 28806 4246 28858
rect 4298 28806 4310 28858
rect 4362 28806 4374 28858
rect 4426 28806 4438 28858
rect 4490 28806 4502 28858
rect 4554 28806 10182 28858
rect 10234 28806 10246 28858
rect 10298 28806 10310 28858
rect 10362 28806 10374 28858
rect 10426 28806 10438 28858
rect 10490 28806 10502 28858
rect 10554 28806 16182 28858
rect 16234 28806 16246 28858
rect 16298 28806 16310 28858
rect 16362 28806 16374 28858
rect 16426 28806 16438 28858
rect 16490 28806 16502 28858
rect 16554 28806 22182 28858
rect 22234 28806 22246 28858
rect 22298 28806 22310 28858
rect 22362 28806 22374 28858
rect 22426 28806 22438 28858
rect 22490 28806 22502 28858
rect 22554 28806 28182 28858
rect 28234 28806 28246 28858
rect 28298 28806 28310 28858
rect 28362 28806 28374 28858
rect 28426 28806 28438 28858
rect 28490 28806 28502 28858
rect 28554 28806 31280 28858
rect 1104 28784 31280 28806
rect 7006 28704 7012 28756
rect 7064 28704 7070 28756
rect 8478 28704 8484 28756
rect 8536 28744 8542 28756
rect 8941 28747 8999 28753
rect 8941 28744 8953 28747
rect 8536 28716 8953 28744
rect 8536 28704 8542 28716
rect 8941 28713 8953 28716
rect 8987 28713 8999 28747
rect 8941 28707 8999 28713
rect 10505 28747 10563 28753
rect 10505 28713 10517 28747
rect 10551 28744 10563 28747
rect 10594 28744 10600 28756
rect 10551 28716 10600 28744
rect 10551 28713 10563 28716
rect 10505 28707 10563 28713
rect 10594 28704 10600 28716
rect 10652 28704 10658 28756
rect 12989 28747 13047 28753
rect 12989 28713 13001 28747
rect 13035 28744 13047 28747
rect 13170 28744 13176 28756
rect 13035 28716 13176 28744
rect 13035 28713 13047 28716
rect 12989 28707 13047 28713
rect 13170 28704 13176 28716
rect 13228 28704 13234 28756
rect 15473 28747 15531 28753
rect 15473 28713 15485 28747
rect 15519 28744 15531 28747
rect 15565 28747 15623 28753
rect 15565 28744 15577 28747
rect 15519 28716 15577 28744
rect 15519 28713 15531 28716
rect 15473 28707 15531 28713
rect 15565 28713 15577 28716
rect 15611 28713 15623 28747
rect 15565 28707 15623 28713
rect 18785 28747 18843 28753
rect 18785 28713 18797 28747
rect 18831 28744 18843 28747
rect 19794 28744 19800 28756
rect 18831 28716 19800 28744
rect 18831 28713 18843 28716
rect 18785 28707 18843 28713
rect 19794 28704 19800 28716
rect 19852 28704 19858 28756
rect 20809 28747 20867 28753
rect 20809 28713 20821 28747
rect 20855 28744 20867 28747
rect 20990 28744 20996 28756
rect 20855 28716 20996 28744
rect 20855 28713 20867 28716
rect 20809 28707 20867 28713
rect 20990 28704 20996 28716
rect 21048 28704 21054 28756
rect 6917 28679 6975 28685
rect 6917 28645 6929 28679
rect 6963 28676 6975 28679
rect 6963 28648 8432 28676
rect 6963 28645 6975 28648
rect 6917 28639 6975 28645
rect 8404 28620 8432 28648
rect 11330 28636 11336 28688
rect 11388 28676 11394 28688
rect 12621 28679 12679 28685
rect 11388 28648 12480 28676
rect 11388 28636 11394 28648
rect 7374 28608 7380 28620
rect 6564 28580 7380 28608
rect 5537 28543 5595 28549
rect 5537 28509 5549 28543
rect 5583 28540 5595 28543
rect 6564 28540 6592 28580
rect 7374 28568 7380 28580
rect 7432 28568 7438 28620
rect 7466 28568 7472 28620
rect 7524 28608 7530 28620
rect 7561 28611 7619 28617
rect 7561 28608 7573 28611
rect 7524 28580 7573 28608
rect 7524 28568 7530 28580
rect 7561 28577 7573 28580
rect 7607 28577 7619 28611
rect 7561 28571 7619 28577
rect 8386 28568 8392 28620
rect 8444 28568 8450 28620
rect 9585 28611 9643 28617
rect 9585 28577 9597 28611
rect 9631 28608 9643 28611
rect 9950 28608 9956 28620
rect 9631 28580 9956 28608
rect 9631 28577 9643 28580
rect 9585 28571 9643 28577
rect 9950 28568 9956 28580
rect 10008 28608 10014 28620
rect 12158 28608 12164 28620
rect 10008 28580 12164 28608
rect 10008 28568 10014 28580
rect 12158 28568 12164 28580
rect 12216 28568 12222 28620
rect 5583 28512 6592 28540
rect 9309 28543 9367 28549
rect 5583 28509 5595 28512
rect 5537 28503 5595 28509
rect 9309 28509 9321 28543
rect 9355 28540 9367 28543
rect 9398 28540 9404 28552
rect 9355 28512 9404 28540
rect 9355 28509 9367 28512
rect 9309 28503 9367 28509
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28540 10747 28543
rect 11514 28540 11520 28552
rect 10735 28512 11520 28540
rect 10735 28509 10747 28512
rect 10689 28503 10747 28509
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 12066 28500 12072 28552
rect 12124 28500 12130 28552
rect 12342 28500 12348 28552
rect 12400 28500 12406 28552
rect 12452 28549 12480 28648
rect 12621 28645 12633 28679
rect 12667 28676 12679 28679
rect 19812 28676 19840 28704
rect 12667 28648 15884 28676
rect 19812 28648 20760 28676
rect 12667 28645 12679 28648
rect 12621 28639 12679 28645
rect 13170 28608 13176 28620
rect 12728 28580 13176 28608
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28509 12495 28543
rect 12437 28503 12495 28509
rect 5804 28475 5862 28481
rect 5804 28441 5816 28475
rect 5850 28472 5862 28475
rect 6362 28472 6368 28484
rect 5850 28444 6368 28472
rect 5850 28441 5862 28444
rect 5804 28435 5862 28441
rect 6362 28432 6368 28444
rect 6420 28432 6426 28484
rect 8478 28472 8484 28484
rect 7392 28444 8484 28472
rect 7392 28413 7420 28444
rect 8478 28432 8484 28444
rect 8536 28472 8542 28484
rect 11974 28472 11980 28484
rect 8536 28444 11980 28472
rect 8536 28432 8542 28444
rect 11974 28432 11980 28444
rect 12032 28432 12038 28484
rect 12158 28432 12164 28484
rect 12216 28472 12222 28484
rect 12253 28475 12311 28481
rect 12253 28472 12265 28475
rect 12216 28444 12265 28472
rect 12216 28432 12222 28444
rect 12253 28441 12265 28444
rect 12299 28441 12311 28475
rect 12728 28472 12756 28580
rect 13170 28568 13176 28580
rect 13228 28608 13234 28620
rect 13541 28611 13599 28617
rect 13541 28608 13553 28611
rect 13228 28580 13553 28608
rect 13228 28568 13234 28580
rect 13541 28577 13553 28580
rect 13587 28577 13599 28611
rect 13541 28571 13599 28577
rect 13725 28611 13783 28617
rect 13725 28577 13737 28611
rect 13771 28577 13783 28611
rect 13725 28571 13783 28577
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28540 12863 28543
rect 13740 28540 13768 28571
rect 14458 28568 14464 28620
rect 14516 28608 14522 28620
rect 14645 28611 14703 28617
rect 14645 28608 14657 28611
rect 14516 28580 14657 28608
rect 14516 28568 14522 28580
rect 14645 28577 14657 28580
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 14921 28543 14979 28549
rect 12851 28512 13124 28540
rect 13740 28512 14596 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 12253 28435 12311 28441
rect 12406 28444 12756 28472
rect 7377 28407 7435 28413
rect 7377 28373 7389 28407
rect 7423 28373 7435 28407
rect 7377 28367 7435 28373
rect 7469 28407 7527 28413
rect 7469 28373 7481 28407
rect 7515 28404 7527 28407
rect 7837 28407 7895 28413
rect 7837 28404 7849 28407
rect 7515 28376 7849 28404
rect 7515 28373 7527 28376
rect 7469 28367 7527 28373
rect 7837 28373 7849 28376
rect 7883 28373 7895 28407
rect 7837 28367 7895 28373
rect 8294 28364 8300 28416
rect 8352 28404 8358 28416
rect 9401 28407 9459 28413
rect 9401 28404 9413 28407
rect 8352 28376 9413 28404
rect 8352 28364 8358 28376
rect 9401 28373 9413 28376
rect 9447 28404 9459 28407
rect 12406 28404 12434 28444
rect 13096 28413 13124 28512
rect 13449 28475 13507 28481
rect 13449 28441 13461 28475
rect 13495 28472 13507 28475
rect 14093 28475 14151 28481
rect 14093 28472 14105 28475
rect 13495 28444 14105 28472
rect 13495 28441 13507 28444
rect 13449 28435 13507 28441
rect 14093 28441 14105 28444
rect 14139 28441 14151 28475
rect 14093 28435 14151 28441
rect 14568 28416 14596 28512
rect 14921 28509 14933 28543
rect 14967 28540 14979 28543
rect 15010 28540 15016 28552
rect 14967 28512 15016 28540
rect 14967 28509 14979 28512
rect 14921 28503 14979 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 15102 28500 15108 28552
rect 15160 28500 15166 28552
rect 15194 28500 15200 28552
rect 15252 28500 15258 28552
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 15378 28540 15384 28552
rect 15335 28512 15384 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15378 28500 15384 28512
rect 15436 28540 15442 28552
rect 15436 28512 15700 28540
rect 15436 28500 15442 28512
rect 15562 28432 15568 28484
rect 15620 28432 15626 28484
rect 15672 28472 15700 28512
rect 15746 28500 15752 28552
rect 15804 28500 15810 28552
rect 15856 28549 15884 28648
rect 15948 28580 17540 28608
rect 15841 28543 15899 28549
rect 15841 28509 15853 28543
rect 15887 28509 15899 28543
rect 15841 28503 15899 28509
rect 15948 28472 15976 28580
rect 17310 28500 17316 28552
rect 17368 28540 17374 28552
rect 17405 28543 17463 28549
rect 17405 28540 17417 28543
rect 17368 28512 17417 28540
rect 17368 28500 17374 28512
rect 17405 28509 17417 28512
rect 17451 28509 17463 28543
rect 17512 28540 17540 28580
rect 18874 28568 18880 28620
rect 18932 28608 18938 28620
rect 20732 28617 20760 28648
rect 19797 28611 19855 28617
rect 19797 28608 19809 28611
rect 18932 28580 19809 28608
rect 18932 28568 18938 28580
rect 19797 28577 19809 28580
rect 19843 28577 19855 28611
rect 19797 28571 19855 28577
rect 20717 28611 20775 28617
rect 20717 28577 20729 28611
rect 20763 28577 20775 28611
rect 20717 28571 20775 28577
rect 20898 28568 20904 28620
rect 20956 28608 20962 28620
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 20956 28580 21373 28608
rect 20956 28568 20962 28580
rect 21361 28577 21373 28580
rect 21407 28577 21419 28611
rect 21361 28571 21419 28577
rect 20346 28540 20352 28552
rect 17512 28512 20352 28540
rect 17405 28503 17463 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28540 21235 28543
rect 21818 28540 21824 28552
rect 21223 28512 21824 28540
rect 21223 28509 21235 28512
rect 21177 28503 21235 28509
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 15672 28444 15976 28472
rect 17494 28432 17500 28484
rect 17552 28472 17558 28484
rect 17650 28475 17708 28481
rect 17650 28472 17662 28475
rect 17552 28444 17662 28472
rect 17552 28432 17558 28444
rect 17650 28441 17662 28444
rect 17696 28441 17708 28475
rect 17650 28435 17708 28441
rect 19613 28475 19671 28481
rect 19613 28441 19625 28475
rect 19659 28472 19671 28475
rect 20073 28475 20131 28481
rect 20073 28472 20085 28475
rect 19659 28444 20085 28472
rect 19659 28441 19671 28444
rect 19613 28435 19671 28441
rect 20073 28441 20085 28444
rect 20119 28441 20131 28475
rect 20073 28435 20131 28441
rect 9447 28376 12434 28404
rect 13081 28407 13139 28413
rect 9447 28373 9459 28376
rect 9401 28367 9459 28373
rect 13081 28373 13093 28407
rect 13127 28373 13139 28407
rect 13081 28367 13139 28373
rect 14550 28364 14556 28416
rect 14608 28364 14614 28416
rect 15378 28364 15384 28416
rect 15436 28404 15442 28416
rect 16025 28407 16083 28413
rect 16025 28404 16037 28407
rect 15436 28376 16037 28404
rect 15436 28364 15442 28376
rect 16025 28373 16037 28376
rect 16071 28373 16083 28407
rect 16025 28367 16083 28373
rect 19242 28364 19248 28416
rect 19300 28364 19306 28416
rect 19702 28364 19708 28416
rect 19760 28364 19766 28416
rect 21269 28407 21327 28413
rect 21269 28373 21281 28407
rect 21315 28404 21327 28407
rect 22094 28404 22100 28416
rect 21315 28376 22100 28404
rect 21315 28373 21327 28376
rect 21269 28367 21327 28373
rect 22094 28364 22100 28376
rect 22152 28364 22158 28416
rect 1104 28314 31280 28336
rect 1104 28262 4922 28314
rect 4974 28262 4986 28314
rect 5038 28262 5050 28314
rect 5102 28262 5114 28314
rect 5166 28262 5178 28314
rect 5230 28262 5242 28314
rect 5294 28262 10922 28314
rect 10974 28262 10986 28314
rect 11038 28262 11050 28314
rect 11102 28262 11114 28314
rect 11166 28262 11178 28314
rect 11230 28262 11242 28314
rect 11294 28262 16922 28314
rect 16974 28262 16986 28314
rect 17038 28262 17050 28314
rect 17102 28262 17114 28314
rect 17166 28262 17178 28314
rect 17230 28262 17242 28314
rect 17294 28262 22922 28314
rect 22974 28262 22986 28314
rect 23038 28262 23050 28314
rect 23102 28262 23114 28314
rect 23166 28262 23178 28314
rect 23230 28262 23242 28314
rect 23294 28262 28922 28314
rect 28974 28262 28986 28314
rect 29038 28262 29050 28314
rect 29102 28262 29114 28314
rect 29166 28262 29178 28314
rect 29230 28262 29242 28314
rect 29294 28262 31280 28314
rect 1104 28240 31280 28262
rect 5534 28160 5540 28212
rect 5592 28200 5598 28212
rect 5721 28203 5779 28209
rect 5721 28200 5733 28203
rect 5592 28172 5733 28200
rect 5592 28160 5598 28172
rect 5721 28169 5733 28172
rect 5767 28169 5779 28203
rect 5721 28163 5779 28169
rect 5813 28203 5871 28209
rect 5813 28169 5825 28203
rect 5859 28200 5871 28203
rect 6362 28200 6368 28212
rect 5859 28172 6368 28200
rect 5859 28169 5871 28172
rect 5813 28163 5871 28169
rect 6362 28160 6368 28172
rect 6420 28160 6426 28212
rect 6546 28160 6552 28212
rect 6604 28200 6610 28212
rect 8294 28200 8300 28212
rect 6604 28172 8300 28200
rect 6604 28160 6610 28172
rect 8294 28160 8300 28172
rect 8352 28160 8358 28212
rect 8386 28160 8392 28212
rect 8444 28160 8450 28212
rect 9125 28203 9183 28209
rect 9125 28169 9137 28203
rect 9171 28200 9183 28203
rect 15562 28200 15568 28212
rect 9171 28172 15568 28200
rect 9171 28169 9183 28172
rect 9125 28163 9183 28169
rect 15562 28160 15568 28172
rect 15620 28160 15626 28212
rect 17405 28203 17463 28209
rect 17405 28169 17417 28203
rect 17451 28200 17463 28203
rect 17494 28200 17500 28212
rect 17451 28172 17500 28200
rect 17451 28169 17463 28172
rect 17405 28163 17463 28169
rect 17494 28160 17500 28172
rect 17552 28160 17558 28212
rect 19242 28200 19248 28212
rect 17604 28172 19248 28200
rect 8404 28132 8432 28160
rect 8849 28135 8907 28141
rect 8849 28132 8861 28135
rect 3896 28104 7420 28132
rect 8404 28104 8861 28132
rect 3896 28073 3924 28104
rect 3881 28067 3939 28073
rect 3881 28033 3893 28067
rect 3927 28033 3939 28067
rect 3881 28027 3939 28033
rect 4148 28067 4206 28073
rect 4148 28033 4160 28067
rect 4194 28064 4206 28067
rect 4614 28064 4620 28076
rect 4194 28036 4620 28064
rect 4194 28033 4206 28036
rect 4148 28027 4206 28033
rect 4614 28024 4620 28036
rect 4672 28024 4678 28076
rect 6380 28073 6408 28104
rect 7392 28076 7420 28104
rect 8849 28101 8861 28104
rect 8895 28101 8907 28135
rect 8849 28095 8907 28101
rect 12805 28135 12863 28141
rect 12805 28101 12817 28135
rect 12851 28132 12863 28135
rect 13630 28132 13636 28144
rect 12851 28104 13636 28132
rect 12851 28101 12863 28104
rect 12805 28095 12863 28101
rect 13630 28092 13636 28104
rect 13688 28092 13694 28144
rect 6365 28067 6423 28073
rect 6365 28033 6377 28067
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 6454 28024 6460 28076
rect 6512 28064 6518 28076
rect 6621 28067 6679 28073
rect 6621 28064 6633 28067
rect 6512 28036 6633 28064
rect 6512 28024 6518 28036
rect 6621 28033 6633 28036
rect 6667 28033 6679 28067
rect 6621 28027 6679 28033
rect 7374 28024 7380 28076
rect 7432 28024 7438 28076
rect 7650 28024 7656 28076
rect 7708 28064 7714 28076
rect 7708 28036 8524 28064
rect 7708 28024 7714 28036
rect 5994 27956 6000 28008
rect 6052 27956 6058 28008
rect 8389 27999 8447 28005
rect 8389 27965 8401 27999
rect 8435 27965 8447 27999
rect 8496 27996 8524 28036
rect 8570 28024 8576 28076
rect 8628 28024 8634 28076
rect 8754 28024 8760 28076
rect 8812 28024 8818 28076
rect 8941 28067 8999 28073
rect 8941 28033 8953 28067
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 8956 27996 8984 28027
rect 9122 28024 9128 28076
rect 9180 28064 9186 28076
rect 10689 28067 10747 28073
rect 10689 28064 10701 28067
rect 9180 28036 10701 28064
rect 9180 28024 9186 28036
rect 10689 28033 10701 28036
rect 10735 28033 10747 28067
rect 10965 28067 11023 28073
rect 10965 28064 10977 28067
rect 10689 28027 10747 28033
rect 10796 28036 10977 28064
rect 10796 27996 10824 28036
rect 10965 28033 10977 28036
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 12621 28067 12679 28073
rect 12621 28033 12633 28067
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28064 12955 28067
rect 13722 28064 13728 28076
rect 12943 28036 13728 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 8496 27968 8984 27996
rect 10704 27968 10824 27996
rect 10873 27999 10931 28005
rect 8389 27959 8447 27965
rect 5261 27931 5319 27937
rect 5261 27897 5273 27931
rect 5307 27928 5319 27931
rect 5307 27900 6132 27928
rect 5307 27897 5319 27900
rect 5261 27891 5319 27897
rect 6104 27872 6132 27900
rect 7742 27888 7748 27940
rect 7800 27928 7806 27940
rect 8404 27928 8432 27959
rect 10704 27940 10732 27968
rect 10873 27965 10885 27999
rect 10919 27996 10931 27999
rect 12437 27999 12495 28005
rect 12437 27996 12449 27999
rect 10919 27968 12449 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 12437 27965 12449 27968
rect 12483 27965 12495 27999
rect 12636 27996 12664 28027
rect 13722 28024 13728 28036
rect 13780 28024 13786 28076
rect 17221 28067 17279 28073
rect 17221 28033 17233 28067
rect 17267 28064 17279 28067
rect 17604 28064 17632 28172
rect 19242 28160 19248 28172
rect 19300 28160 19306 28212
rect 22373 28203 22431 28209
rect 22373 28169 22385 28203
rect 22419 28200 22431 28203
rect 22419 28172 23612 28200
rect 22419 28169 22431 28172
rect 22373 28163 22431 28169
rect 17678 28092 17684 28144
rect 17736 28132 17742 28144
rect 17736 28104 17816 28132
rect 17736 28092 17742 28104
rect 17788 28073 17816 28104
rect 22278 28092 22284 28144
rect 22336 28132 22342 28144
rect 23584 28141 23612 28172
rect 23569 28135 23627 28141
rect 22336 28104 23152 28132
rect 22336 28092 22342 28104
rect 17267 28036 17632 28064
rect 17764 28067 17822 28073
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 17764 28033 17776 28067
rect 17810 28033 17822 28067
rect 17764 28027 17822 28033
rect 21634 28024 21640 28076
rect 21692 28064 21698 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21692 28036 21833 28064
rect 21692 28024 21698 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22097 28067 22155 28073
rect 22097 28033 22109 28067
rect 22143 28033 22155 28067
rect 22097 28027 22155 28033
rect 22189 28067 22247 28073
rect 22189 28033 22201 28067
rect 22235 28064 22247 28067
rect 22462 28064 22468 28076
rect 22235 28036 22468 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 13538 27996 13544 28008
rect 12636 27968 13544 27996
rect 12437 27959 12495 27965
rect 13538 27956 13544 27968
rect 13596 27956 13602 28008
rect 17310 27956 17316 28008
rect 17368 27996 17374 28008
rect 17497 27999 17555 28005
rect 17497 27996 17509 27999
rect 17368 27968 17509 27996
rect 17368 27956 17374 27968
rect 17497 27965 17509 27968
rect 17543 27965 17555 27999
rect 22020 27996 22048 28027
rect 17497 27959 17555 27965
rect 21836 27968 22048 27996
rect 22112 27996 22140 28027
rect 22462 28024 22468 28036
rect 22520 28024 22526 28076
rect 22646 28024 22652 28076
rect 22704 28024 22710 28076
rect 22922 28024 22928 28076
rect 22980 28024 22986 28076
rect 22664 27996 22692 28024
rect 22112 27968 22692 27996
rect 23017 27999 23075 28005
rect 21836 27940 21864 27968
rect 23017 27965 23029 27999
rect 23063 27965 23075 27999
rect 23124 27996 23152 28104
rect 23569 28101 23581 28135
rect 23615 28101 23627 28135
rect 23569 28095 23627 28101
rect 23201 28067 23259 28073
rect 23201 28033 23213 28067
rect 23247 28064 23259 28067
rect 23382 28064 23388 28076
rect 23247 28036 23388 28064
rect 23247 28033 23259 28036
rect 23201 28027 23259 28033
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28064 23903 28067
rect 24026 28064 24032 28076
rect 23891 28036 24032 28064
rect 23891 28033 23903 28036
rect 23845 28027 23903 28033
rect 24026 28024 24032 28036
rect 24084 28024 24090 28076
rect 23124 27968 23612 27996
rect 23017 27959 23075 27965
rect 7800 27900 8432 27928
rect 7800 27888 7806 27900
rect 10686 27888 10692 27940
rect 10744 27888 10750 27940
rect 18877 27931 18935 27937
rect 10980 27900 11652 27928
rect 5350 27820 5356 27872
rect 5408 27820 5414 27872
rect 6086 27820 6092 27872
rect 6144 27820 6150 27872
rect 7834 27820 7840 27872
rect 7892 27820 7898 27872
rect 10980 27869 11008 27900
rect 11624 27872 11652 27900
rect 18877 27897 18889 27931
rect 18923 27928 18935 27931
rect 19334 27928 19340 27940
rect 18923 27900 19340 27928
rect 18923 27897 18935 27900
rect 18877 27891 18935 27897
rect 19334 27888 19340 27900
rect 19392 27888 19398 27940
rect 21818 27888 21824 27940
rect 21876 27888 21882 27940
rect 23032 27928 23060 27959
rect 23474 27928 23480 27940
rect 22066 27900 22968 27928
rect 23032 27900 23480 27928
rect 10965 27863 11023 27869
rect 10965 27829 10977 27863
rect 11011 27829 11023 27863
rect 10965 27823 11023 27829
rect 11146 27820 11152 27872
rect 11204 27820 11210 27872
rect 11606 27820 11612 27872
rect 11664 27820 11670 27872
rect 20714 27820 20720 27872
rect 20772 27860 20778 27872
rect 22066 27860 22094 27900
rect 22940 27869 22968 27900
rect 23474 27888 23480 27900
rect 23532 27888 23538 27940
rect 20772 27832 22094 27860
rect 22925 27863 22983 27869
rect 20772 27820 20778 27832
rect 22925 27829 22937 27863
rect 22971 27829 22983 27863
rect 22925 27823 22983 27829
rect 23014 27820 23020 27872
rect 23072 27860 23078 27872
rect 23584 27869 23612 27968
rect 23750 27956 23756 28008
rect 23808 27956 23814 28008
rect 23385 27863 23443 27869
rect 23385 27860 23397 27863
rect 23072 27832 23397 27860
rect 23072 27820 23078 27832
rect 23385 27829 23397 27832
rect 23431 27829 23443 27863
rect 23385 27823 23443 27829
rect 23569 27863 23627 27869
rect 23569 27829 23581 27863
rect 23615 27829 23627 27863
rect 23569 27823 23627 27829
rect 24026 27820 24032 27872
rect 24084 27820 24090 27872
rect 1104 27770 31280 27792
rect 1104 27718 4182 27770
rect 4234 27718 4246 27770
rect 4298 27718 4310 27770
rect 4362 27718 4374 27770
rect 4426 27718 4438 27770
rect 4490 27718 4502 27770
rect 4554 27718 10182 27770
rect 10234 27718 10246 27770
rect 10298 27718 10310 27770
rect 10362 27718 10374 27770
rect 10426 27718 10438 27770
rect 10490 27718 10502 27770
rect 10554 27718 16182 27770
rect 16234 27718 16246 27770
rect 16298 27718 16310 27770
rect 16362 27718 16374 27770
rect 16426 27718 16438 27770
rect 16490 27718 16502 27770
rect 16554 27718 22182 27770
rect 22234 27718 22246 27770
rect 22298 27718 22310 27770
rect 22362 27718 22374 27770
rect 22426 27718 22438 27770
rect 22490 27718 22502 27770
rect 22554 27718 28182 27770
rect 28234 27718 28246 27770
rect 28298 27718 28310 27770
rect 28362 27718 28374 27770
rect 28426 27718 28438 27770
rect 28490 27718 28502 27770
rect 28554 27718 31280 27770
rect 1104 27696 31280 27718
rect 4249 27659 4307 27665
rect 4249 27625 4261 27659
rect 4295 27656 4307 27659
rect 4614 27656 4620 27668
rect 4295 27628 4620 27656
rect 4295 27625 4307 27628
rect 4249 27619 4307 27625
rect 4614 27616 4620 27628
rect 4672 27616 4678 27668
rect 6089 27659 6147 27665
rect 6089 27625 6101 27659
rect 6135 27656 6147 27659
rect 6454 27656 6460 27668
rect 6135 27628 6460 27656
rect 6135 27625 6147 27628
rect 6089 27619 6147 27625
rect 6454 27616 6460 27628
rect 6512 27616 6518 27668
rect 7190 27616 7196 27668
rect 7248 27656 7254 27668
rect 8754 27656 8760 27668
rect 7248 27628 8760 27656
rect 7248 27616 7254 27628
rect 8754 27616 8760 27628
rect 8812 27616 8818 27668
rect 9122 27616 9128 27668
rect 9180 27616 9186 27668
rect 13630 27616 13636 27668
rect 13688 27616 13694 27668
rect 15746 27616 15752 27668
rect 15804 27656 15810 27668
rect 16393 27659 16451 27665
rect 16393 27656 16405 27659
rect 15804 27628 16405 27656
rect 15804 27616 15810 27628
rect 16393 27625 16405 27628
rect 16439 27625 16451 27659
rect 16393 27619 16451 27625
rect 22002 27616 22008 27668
rect 22060 27616 22066 27668
rect 22922 27616 22928 27668
rect 22980 27656 22986 27668
rect 23385 27659 23443 27665
rect 23385 27656 23397 27659
rect 22980 27628 23397 27656
rect 22980 27616 22986 27628
rect 23385 27625 23397 27628
rect 23431 27625 23443 27659
rect 23385 27619 23443 27625
rect 6181 27591 6239 27597
rect 6181 27557 6193 27591
rect 6227 27557 6239 27591
rect 7466 27588 7472 27600
rect 6181 27551 6239 27557
rect 6840 27560 7472 27588
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27452 4491 27455
rect 5350 27452 5356 27464
rect 4479 27424 5356 27452
rect 4479 27421 4491 27424
rect 4433 27415 4491 27421
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 5905 27455 5963 27461
rect 5905 27421 5917 27455
rect 5951 27452 5963 27455
rect 6196 27452 6224 27551
rect 6840 27529 6868 27560
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 7561 27591 7619 27597
rect 7561 27557 7573 27591
rect 7607 27588 7619 27591
rect 9140 27588 9168 27616
rect 7607 27560 9168 27588
rect 7607 27557 7619 27560
rect 7561 27551 7619 27557
rect 6825 27523 6883 27529
rect 6825 27489 6837 27523
rect 6871 27489 6883 27523
rect 7834 27520 7840 27532
rect 6825 27483 6883 27489
rect 6932 27492 7840 27520
rect 5951 27424 6224 27452
rect 6641 27455 6699 27461
rect 5951 27421 5963 27424
rect 5905 27415 5963 27421
rect 6641 27421 6653 27455
rect 6687 27452 6699 27455
rect 6932 27452 6960 27492
rect 7834 27480 7840 27492
rect 7892 27480 7898 27532
rect 13648 27520 13676 27616
rect 13722 27548 13728 27600
rect 13780 27588 13786 27600
rect 13780 27560 15240 27588
rect 13780 27548 13786 27560
rect 14645 27523 14703 27529
rect 14645 27520 14657 27523
rect 13648 27492 14657 27520
rect 14645 27489 14657 27492
rect 14691 27489 14703 27523
rect 15212 27520 15240 27560
rect 16574 27548 16580 27600
rect 16632 27588 16638 27600
rect 22370 27588 22376 27600
rect 16632 27560 22376 27588
rect 16632 27548 16638 27560
rect 22370 27548 22376 27560
rect 22428 27548 22434 27600
rect 22572 27560 24992 27588
rect 15212 27492 16896 27520
rect 14645 27483 14703 27489
rect 6687 27424 6960 27452
rect 7009 27455 7067 27461
rect 6687 27421 6699 27424
rect 6641 27415 6699 27421
rect 7009 27421 7021 27455
rect 7055 27421 7067 27455
rect 7009 27415 7067 27421
rect 6086 27344 6092 27396
rect 6144 27384 6150 27396
rect 7024 27384 7052 27415
rect 7190 27412 7196 27464
rect 7248 27412 7254 27464
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 7650 27452 7656 27464
rect 7423 27424 7656 27452
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 7650 27412 7656 27424
rect 7708 27412 7714 27464
rect 7742 27412 7748 27464
rect 7800 27412 7806 27464
rect 11974 27412 11980 27464
rect 12032 27412 12038 27464
rect 12253 27455 12311 27461
rect 12253 27421 12265 27455
rect 12299 27452 12311 27455
rect 12342 27452 12348 27464
rect 12299 27424 12348 27452
rect 12299 27421 12311 27424
rect 12253 27415 12311 27421
rect 12342 27412 12348 27424
rect 12400 27412 12406 27464
rect 15746 27412 15752 27464
rect 15804 27452 15810 27464
rect 15804 27424 16436 27452
rect 15804 27412 15810 27424
rect 6144 27356 7052 27384
rect 7285 27387 7343 27393
rect 6144 27344 6150 27356
rect 7285 27353 7297 27387
rect 7331 27384 7343 27387
rect 7760 27384 7788 27412
rect 12498 27387 12556 27393
rect 12498 27384 12510 27387
rect 7331 27356 7788 27384
rect 12406 27356 12510 27384
rect 7331 27353 7343 27356
rect 7285 27347 7343 27353
rect 6546 27276 6552 27328
rect 6604 27276 6610 27328
rect 12161 27319 12219 27325
rect 12161 27285 12173 27319
rect 12207 27316 12219 27319
rect 12406 27316 12434 27356
rect 12498 27353 12510 27356
rect 12544 27353 12556 27387
rect 12498 27347 12556 27353
rect 12207 27288 12434 27316
rect 12207 27285 12219 27288
rect 12161 27279 12219 27285
rect 14090 27276 14096 27328
rect 14148 27276 14154 27328
rect 16022 27276 16028 27328
rect 16080 27316 16086 27328
rect 16301 27319 16359 27325
rect 16301 27316 16313 27319
rect 16080 27288 16313 27316
rect 16080 27276 16086 27288
rect 16301 27285 16313 27288
rect 16347 27285 16359 27319
rect 16408 27316 16436 27424
rect 16574 27412 16580 27464
rect 16632 27412 16638 27464
rect 16868 27461 16896 27492
rect 20990 27480 20996 27532
rect 21048 27520 21054 27532
rect 21361 27523 21419 27529
rect 21361 27520 21373 27523
rect 21048 27492 21373 27520
rect 21048 27480 21054 27492
rect 21361 27489 21373 27492
rect 21407 27489 21419 27523
rect 22572 27520 22600 27560
rect 21361 27483 21419 27489
rect 21468 27492 22600 27520
rect 16853 27455 16911 27461
rect 16853 27421 16865 27455
rect 16899 27421 16911 27455
rect 16853 27415 16911 27421
rect 17129 27455 17187 27461
rect 17129 27421 17141 27455
rect 17175 27421 17187 27455
rect 17129 27415 17187 27421
rect 16666 27344 16672 27396
rect 16724 27384 16730 27396
rect 17144 27384 17172 27415
rect 19426 27412 19432 27464
rect 19484 27452 19490 27464
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 19484 27424 20821 27452
rect 19484 27412 19490 27424
rect 20809 27421 20821 27424
rect 20855 27452 20867 27455
rect 21468 27452 21496 27492
rect 22646 27480 22652 27532
rect 22704 27520 22710 27532
rect 22741 27523 22799 27529
rect 22741 27520 22753 27523
rect 22704 27492 22753 27520
rect 22704 27480 22710 27492
rect 22741 27489 22753 27492
rect 22787 27489 22799 27523
rect 22922 27520 22928 27532
rect 22741 27483 22799 27489
rect 22848 27492 22928 27520
rect 20855 27424 21496 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21542 27412 21548 27464
rect 21600 27412 21606 27464
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 22848 27461 22876 27492
rect 22922 27480 22928 27492
rect 22980 27480 22986 27532
rect 24854 27480 24860 27532
rect 24912 27480 24918 27532
rect 24964 27464 24992 27560
rect 22833 27455 22891 27461
rect 21968 27424 22416 27452
rect 21968 27412 21974 27424
rect 20901 27387 20959 27393
rect 16724 27356 17172 27384
rect 19720 27356 20576 27384
rect 16724 27344 16730 27356
rect 19720 27328 19748 27356
rect 16761 27319 16819 27325
rect 16761 27316 16773 27319
rect 16408 27288 16773 27316
rect 16301 27279 16359 27285
rect 16761 27285 16773 27288
rect 16807 27285 16819 27319
rect 16761 27279 16819 27285
rect 16850 27276 16856 27328
rect 16908 27316 16914 27328
rect 16945 27319 17003 27325
rect 16945 27316 16957 27319
rect 16908 27288 16957 27316
rect 16908 27276 16914 27288
rect 16945 27285 16957 27288
rect 16991 27285 17003 27319
rect 16945 27279 17003 27285
rect 19702 27276 19708 27328
rect 19760 27276 19766 27328
rect 20438 27276 20444 27328
rect 20496 27276 20502 27328
rect 20548 27316 20576 27356
rect 20901 27353 20913 27387
rect 20947 27384 20959 27387
rect 22097 27387 22155 27393
rect 22097 27384 22109 27387
rect 20947 27356 22109 27384
rect 20947 27353 20959 27356
rect 20901 27347 20959 27353
rect 22097 27353 22109 27356
rect 22143 27353 22155 27387
rect 22388 27384 22416 27424
rect 22833 27421 22845 27455
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 23201 27455 23259 27461
rect 23201 27421 23213 27455
rect 23247 27452 23259 27455
rect 23382 27452 23388 27464
rect 23247 27424 23388 27452
rect 23247 27421 23259 27424
rect 23201 27415 23259 27421
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 24946 27412 24952 27464
rect 25004 27452 25010 27464
rect 25041 27455 25099 27461
rect 25041 27452 25053 27455
rect 25004 27424 25053 27452
rect 25004 27412 25010 27424
rect 25041 27421 25053 27424
rect 25087 27452 25099 27455
rect 25087 27424 25728 27452
rect 25087 27421 25099 27424
rect 25041 27415 25099 27421
rect 23017 27387 23075 27393
rect 23017 27384 23029 27387
rect 22388 27356 23029 27384
rect 22097 27347 22155 27353
rect 23017 27353 23029 27356
rect 23063 27353 23075 27387
rect 23017 27347 23075 27353
rect 23109 27387 23167 27393
rect 23109 27353 23121 27387
rect 23155 27353 23167 27387
rect 23109 27347 23167 27353
rect 25133 27387 25191 27393
rect 25133 27353 25145 27387
rect 25179 27384 25191 27387
rect 25593 27387 25651 27393
rect 25593 27384 25605 27387
rect 25179 27356 25605 27384
rect 25179 27353 25191 27356
rect 25133 27347 25191 27353
rect 25593 27353 25605 27356
rect 25639 27353 25651 27387
rect 25700 27384 25728 27424
rect 26142 27412 26148 27464
rect 26200 27412 26206 27464
rect 25700 27356 26648 27384
rect 25593 27347 25651 27353
rect 21637 27319 21695 27325
rect 21637 27316 21649 27319
rect 20548 27288 21649 27316
rect 21637 27285 21649 27288
rect 21683 27316 21695 27319
rect 22462 27316 22468 27328
rect 21683 27288 22468 27316
rect 21683 27285 21695 27288
rect 21637 27279 21695 27285
rect 22462 27276 22468 27288
rect 22520 27276 22526 27328
rect 22554 27276 22560 27328
rect 22612 27316 22618 27328
rect 23124 27316 23152 27347
rect 22612 27288 23152 27316
rect 25501 27319 25559 27325
rect 22612 27276 22618 27288
rect 25501 27285 25513 27319
rect 25547 27316 25559 27319
rect 26326 27316 26332 27328
rect 25547 27288 26332 27316
rect 25547 27285 25559 27288
rect 25501 27279 25559 27285
rect 26326 27276 26332 27288
rect 26384 27276 26390 27328
rect 26620 27325 26648 27356
rect 26694 27344 26700 27396
rect 26752 27384 26758 27396
rect 27338 27384 27344 27396
rect 26752 27356 27344 27384
rect 26752 27344 26758 27356
rect 27338 27344 27344 27356
rect 27396 27344 27402 27396
rect 26605 27319 26663 27325
rect 26605 27285 26617 27319
rect 26651 27316 26663 27319
rect 27246 27316 27252 27328
rect 26651 27288 27252 27316
rect 26651 27285 26663 27288
rect 26605 27279 26663 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 1104 27226 31280 27248
rect 1104 27174 4922 27226
rect 4974 27174 4986 27226
rect 5038 27174 5050 27226
rect 5102 27174 5114 27226
rect 5166 27174 5178 27226
rect 5230 27174 5242 27226
rect 5294 27174 10922 27226
rect 10974 27174 10986 27226
rect 11038 27174 11050 27226
rect 11102 27174 11114 27226
rect 11166 27174 11178 27226
rect 11230 27174 11242 27226
rect 11294 27174 16922 27226
rect 16974 27174 16986 27226
rect 17038 27174 17050 27226
rect 17102 27174 17114 27226
rect 17166 27174 17178 27226
rect 17230 27174 17242 27226
rect 17294 27174 22922 27226
rect 22974 27174 22986 27226
rect 23038 27174 23050 27226
rect 23102 27174 23114 27226
rect 23166 27174 23178 27226
rect 23230 27174 23242 27226
rect 23294 27174 28922 27226
rect 28974 27174 28986 27226
rect 29038 27174 29050 27226
rect 29102 27174 29114 27226
rect 29166 27174 29178 27226
rect 29230 27174 29242 27226
rect 29294 27174 31280 27226
rect 1104 27152 31280 27174
rect 11974 27072 11980 27124
rect 12032 27112 12038 27124
rect 12713 27115 12771 27121
rect 12713 27112 12725 27115
rect 12032 27084 12725 27112
rect 12032 27072 12038 27084
rect 12713 27081 12725 27084
rect 12759 27081 12771 27115
rect 12713 27075 12771 27081
rect 13081 27115 13139 27121
rect 13081 27081 13093 27115
rect 13127 27112 13139 27115
rect 14090 27112 14096 27124
rect 13127 27084 14096 27112
rect 13127 27081 13139 27084
rect 13081 27075 13139 27081
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 15105 27115 15163 27121
rect 15105 27081 15117 27115
rect 15151 27112 15163 27115
rect 15746 27112 15752 27124
rect 15151 27084 15752 27112
rect 15151 27081 15163 27084
rect 15105 27075 15163 27081
rect 15746 27072 15752 27084
rect 15804 27072 15810 27124
rect 19981 27115 20039 27121
rect 19981 27081 19993 27115
rect 20027 27081 20039 27115
rect 19981 27075 20039 27081
rect 13170 27004 13176 27056
rect 13228 27004 13234 27056
rect 16240 27047 16298 27053
rect 16240 27013 16252 27047
rect 16286 27044 16298 27047
rect 16758 27044 16764 27056
rect 16286 27016 16764 27044
rect 16286 27013 16298 27016
rect 16240 27007 16298 27013
rect 16758 27004 16764 27016
rect 16816 27004 16822 27056
rect 19996 27044 20024 27075
rect 20438 27072 20444 27124
rect 20496 27072 20502 27124
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 21821 27115 21879 27121
rect 21821 27112 21833 27115
rect 21600 27084 21833 27112
rect 21600 27072 21606 27084
rect 21821 27081 21833 27084
rect 21867 27081 21879 27115
rect 21821 27075 21879 27081
rect 22002 27072 22008 27124
rect 22060 27072 22066 27124
rect 22370 27072 22376 27124
rect 22428 27112 22434 27124
rect 22428 27084 23428 27112
rect 22428 27072 22434 27084
rect 20318 27047 20376 27053
rect 20318 27044 20330 27047
rect 19996 27016 20330 27044
rect 20318 27013 20330 27016
rect 20364 27013 20376 27047
rect 20318 27007 20376 27013
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26976 19855 26979
rect 20456 26976 20484 27072
rect 19843 26948 20484 26976
rect 22020 26976 22048 27072
rect 22462 27004 22468 27056
rect 22520 27044 22526 27056
rect 22520 27016 22968 27044
rect 22520 27004 22526 27016
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 22020 26948 22753 26976
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22741 26939 22799 26945
rect 10689 26911 10747 26917
rect 10689 26877 10701 26911
rect 10735 26877 10747 26911
rect 10689 26871 10747 26877
rect 13357 26911 13415 26917
rect 13357 26877 13369 26911
rect 13403 26908 13415 26911
rect 16485 26911 16543 26917
rect 13403 26880 13676 26908
rect 13403 26877 13415 26880
rect 13357 26871 13415 26877
rect 10704 26784 10732 26871
rect 13648 26784 13676 26880
rect 16485 26877 16497 26911
rect 16531 26908 16543 26911
rect 17034 26908 17040 26920
rect 16531 26880 17040 26908
rect 16531 26877 16543 26880
rect 16485 26871 16543 26877
rect 17034 26868 17040 26880
rect 17092 26908 17098 26920
rect 17310 26908 17316 26920
rect 17092 26880 17316 26908
rect 17092 26868 17098 26880
rect 17310 26868 17316 26880
rect 17368 26868 17374 26920
rect 19978 26868 19984 26920
rect 20036 26908 20042 26920
rect 20073 26911 20131 26917
rect 20073 26908 20085 26911
rect 20036 26880 20085 26908
rect 20036 26868 20042 26880
rect 20073 26877 20085 26880
rect 20119 26877 20131 26911
rect 20073 26871 20131 26877
rect 21818 26868 21824 26920
rect 21876 26908 21882 26920
rect 22465 26911 22523 26917
rect 22465 26908 22477 26911
rect 21876 26880 22477 26908
rect 21876 26868 21882 26880
rect 22465 26877 22477 26880
rect 22511 26908 22523 26911
rect 22554 26908 22560 26920
rect 22511 26880 22560 26908
rect 22511 26877 22523 26880
rect 22465 26871 22523 26877
rect 22554 26868 22560 26880
rect 22612 26868 22618 26920
rect 21453 26843 21511 26849
rect 21453 26809 21465 26843
rect 21499 26840 21511 26843
rect 22646 26840 22652 26852
rect 21499 26812 22652 26840
rect 21499 26809 21511 26812
rect 21453 26803 21511 26809
rect 22646 26800 22652 26812
rect 22704 26800 22710 26852
rect 10042 26732 10048 26784
rect 10100 26732 10106 26784
rect 10686 26732 10692 26784
rect 10744 26732 10750 26784
rect 13630 26732 13636 26784
rect 13688 26732 13694 26784
rect 21358 26732 21364 26784
rect 21416 26772 21422 26784
rect 22557 26775 22615 26781
rect 22557 26772 22569 26775
rect 21416 26744 22569 26772
rect 21416 26732 21422 26744
rect 22557 26741 22569 26744
rect 22603 26741 22615 26775
rect 22940 26772 22968 27016
rect 23400 26976 23428 27084
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 23569 27115 23627 27121
rect 23569 27112 23581 27115
rect 23532 27084 23581 27112
rect 23532 27072 23538 27084
rect 23569 27081 23581 27084
rect 23615 27081 23627 27115
rect 23569 27075 23627 27081
rect 23750 27072 23756 27124
rect 23808 27112 23814 27124
rect 24121 27115 24179 27121
rect 24121 27112 24133 27115
rect 23808 27084 24133 27112
rect 23808 27072 23814 27084
rect 24121 27081 24133 27084
rect 24167 27081 24179 27115
rect 24121 27075 24179 27081
rect 24489 27115 24547 27121
rect 24489 27081 24501 27115
rect 24535 27112 24547 27115
rect 24765 27115 24823 27121
rect 24765 27112 24777 27115
rect 24535 27084 24777 27112
rect 24535 27081 24547 27084
rect 24489 27075 24547 27081
rect 24765 27081 24777 27084
rect 24811 27112 24823 27115
rect 26142 27112 26148 27124
rect 24811 27084 26148 27112
rect 24811 27081 24823 27084
rect 24765 27075 24823 27081
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 26237 27115 26295 27121
rect 26237 27081 26249 27115
rect 26283 27081 26295 27115
rect 26237 27075 26295 27081
rect 23937 27047 23995 27053
rect 23937 27013 23949 27047
rect 23983 27044 23995 27047
rect 25774 27044 25780 27056
rect 23983 27016 25780 27044
rect 23983 27013 23995 27016
rect 23937 27007 23995 27013
rect 25774 27004 25780 27016
rect 25832 27004 25838 27056
rect 25900 27047 25958 27053
rect 25900 27013 25912 27047
rect 25946 27044 25958 27047
rect 26252 27044 26280 27075
rect 26326 27072 26332 27124
rect 26384 27072 26390 27124
rect 25946 27016 26280 27044
rect 25946 27013 25958 27016
rect 25900 27007 25958 27013
rect 23753 26979 23811 26985
rect 23753 26976 23765 26979
rect 23400 26948 23765 26976
rect 23753 26945 23765 26948
rect 23799 26945 23811 26979
rect 23753 26939 23811 26945
rect 24029 26979 24087 26985
rect 24029 26945 24041 26979
rect 24075 26976 24087 26979
rect 24305 26980 24363 26985
rect 24394 26980 24400 26988
rect 24305 26979 24400 26980
rect 24075 26948 24256 26976
rect 24075 26945 24087 26948
rect 24029 26939 24087 26945
rect 23768 26840 23796 26939
rect 24228 26920 24256 26948
rect 24305 26945 24317 26979
rect 24351 26952 24400 26979
rect 24351 26945 24363 26952
rect 24305 26939 24363 26945
rect 24394 26936 24400 26952
rect 24452 26936 24458 26988
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 26145 26979 26203 26985
rect 26145 26976 26157 26979
rect 24581 26939 24639 26945
rect 25056 26948 26157 26976
rect 24210 26868 24216 26920
rect 24268 26908 24274 26920
rect 24596 26908 24624 26939
rect 25056 26920 25084 26948
rect 26145 26945 26157 26948
rect 26191 26945 26203 26979
rect 26344 26976 26372 27072
rect 26421 26979 26479 26985
rect 26421 26976 26433 26979
rect 26344 26948 26433 26976
rect 26145 26939 26203 26945
rect 26421 26945 26433 26948
rect 26467 26945 26479 26979
rect 26421 26939 26479 26945
rect 24268 26880 24624 26908
rect 24268 26868 24274 26880
rect 25038 26868 25044 26920
rect 25096 26868 25102 26920
rect 24394 26840 24400 26852
rect 23768 26812 24400 26840
rect 24394 26800 24400 26812
rect 24452 26840 24458 26852
rect 24762 26840 24768 26852
rect 24452 26812 24768 26840
rect 24452 26800 24458 26812
rect 24762 26800 24768 26812
rect 24820 26800 24826 26852
rect 23842 26772 23848 26784
rect 22940 26744 23848 26772
rect 22557 26735 22615 26741
rect 23842 26732 23848 26744
rect 23900 26772 23906 26784
rect 24486 26772 24492 26784
rect 23900 26744 24492 26772
rect 23900 26732 23906 26744
rect 24486 26732 24492 26744
rect 24544 26732 24550 26784
rect 1104 26682 31280 26704
rect 1104 26630 4182 26682
rect 4234 26630 4246 26682
rect 4298 26630 4310 26682
rect 4362 26630 4374 26682
rect 4426 26630 4438 26682
rect 4490 26630 4502 26682
rect 4554 26630 10182 26682
rect 10234 26630 10246 26682
rect 10298 26630 10310 26682
rect 10362 26630 10374 26682
rect 10426 26630 10438 26682
rect 10490 26630 10502 26682
rect 10554 26630 16182 26682
rect 16234 26630 16246 26682
rect 16298 26630 16310 26682
rect 16362 26630 16374 26682
rect 16426 26630 16438 26682
rect 16490 26630 16502 26682
rect 16554 26630 22182 26682
rect 22234 26630 22246 26682
rect 22298 26630 22310 26682
rect 22362 26630 22374 26682
rect 22426 26630 22438 26682
rect 22490 26630 22502 26682
rect 22554 26630 28182 26682
rect 28234 26630 28246 26682
rect 28298 26630 28310 26682
rect 28362 26630 28374 26682
rect 28426 26630 28438 26682
rect 28490 26630 28502 26682
rect 28554 26630 31280 26682
rect 1104 26608 31280 26630
rect 11422 26528 11428 26580
rect 11480 26568 11486 26580
rect 16485 26571 16543 26577
rect 11480 26540 11560 26568
rect 11480 26528 11486 26540
rect 10321 26503 10379 26509
rect 10321 26469 10333 26503
rect 10367 26500 10379 26503
rect 10686 26500 10692 26512
rect 10367 26472 10692 26500
rect 10367 26469 10379 26472
rect 10321 26463 10379 26469
rect 10686 26460 10692 26472
rect 10744 26500 10750 26512
rect 10744 26472 11468 26500
rect 10744 26460 10750 26472
rect 8570 26324 8576 26376
rect 8628 26324 8634 26376
rect 8941 26367 8999 26373
rect 8941 26333 8953 26367
rect 8987 26364 8999 26367
rect 9582 26364 9588 26376
rect 8987 26336 9588 26364
rect 8987 26333 8999 26336
rect 8941 26327 8999 26333
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 10502 26324 10508 26376
rect 10560 26364 10566 26376
rect 11440 26373 11468 26472
rect 11532 26376 11560 26540
rect 16485 26537 16497 26571
rect 16531 26568 16543 26571
rect 16666 26568 16672 26580
rect 16531 26540 16672 26568
rect 16531 26537 16543 26540
rect 16485 26531 16543 26537
rect 16666 26528 16672 26540
rect 16724 26528 16730 26580
rect 18969 26571 19027 26577
rect 18969 26537 18981 26571
rect 19015 26568 19027 26571
rect 19702 26568 19708 26580
rect 19015 26540 19708 26568
rect 19015 26537 19027 26540
rect 18969 26531 19027 26537
rect 19702 26528 19708 26540
rect 19760 26528 19766 26580
rect 21818 26528 21824 26580
rect 21876 26528 21882 26580
rect 25038 26568 25044 26580
rect 22066 26540 25044 26568
rect 13630 26460 13636 26512
rect 13688 26500 13694 26512
rect 15194 26500 15200 26512
rect 13688 26472 15200 26500
rect 13688 26460 13694 26472
rect 13740 26441 13768 26472
rect 15194 26460 15200 26472
rect 15252 26500 15258 26512
rect 20254 26500 20260 26512
rect 15252 26472 20260 26500
rect 15252 26460 15258 26472
rect 13725 26435 13783 26441
rect 13725 26401 13737 26435
rect 13771 26401 13783 26435
rect 13725 26395 13783 26401
rect 15286 26392 15292 26444
rect 15344 26392 15350 26444
rect 15948 26441 15976 26472
rect 20254 26460 20260 26472
rect 20312 26460 20318 26512
rect 15933 26435 15991 26441
rect 15933 26401 15945 26435
rect 15979 26401 15991 26435
rect 15933 26395 15991 26401
rect 16022 26392 16028 26444
rect 16080 26392 16086 26444
rect 17034 26392 17040 26444
rect 17092 26392 17098 26444
rect 11057 26367 11115 26373
rect 11057 26364 11069 26367
rect 10560 26336 11069 26364
rect 10560 26324 10566 26336
rect 11057 26333 11069 26336
rect 11103 26364 11115 26367
rect 11149 26367 11207 26373
rect 11149 26364 11161 26367
rect 11103 26336 11161 26364
rect 11103 26333 11115 26336
rect 11057 26327 11115 26333
rect 11149 26333 11161 26336
rect 11195 26333 11207 26367
rect 11149 26327 11207 26333
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26333 11483 26367
rect 11425 26327 11483 26333
rect 11514 26324 11520 26376
rect 11572 26324 11578 26376
rect 12434 26324 12440 26376
rect 12492 26364 12498 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 12492 26336 13553 26364
rect 12492 26324 12498 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 14642 26324 14648 26376
rect 14700 26324 14706 26376
rect 9186 26299 9244 26305
rect 9186 26296 9198 26299
rect 8772 26268 9198 26296
rect 8772 26237 8800 26268
rect 9186 26265 9198 26268
rect 9232 26265 9244 26299
rect 9186 26259 9244 26265
rect 11333 26299 11391 26305
rect 11333 26265 11345 26299
rect 11379 26296 11391 26299
rect 11790 26296 11796 26308
rect 11379 26268 11796 26296
rect 11379 26265 11391 26268
rect 11333 26259 11391 26265
rect 11790 26256 11796 26268
rect 11848 26296 11854 26308
rect 12158 26296 12164 26308
rect 11848 26268 12164 26296
rect 11848 26256 11854 26268
rect 12158 26256 12164 26268
rect 12216 26256 12222 26308
rect 13449 26299 13507 26305
rect 13449 26265 13461 26299
rect 13495 26296 13507 26299
rect 14093 26299 14151 26305
rect 14093 26296 14105 26299
rect 13495 26268 14105 26296
rect 13495 26265 13507 26268
rect 13449 26259 13507 26265
rect 14093 26265 14105 26268
rect 14139 26265 14151 26299
rect 15304 26296 15332 26392
rect 16040 26364 16068 26392
rect 16117 26367 16175 26373
rect 16117 26364 16129 26367
rect 16040 26336 16129 26364
rect 16117 26333 16129 26336
rect 16163 26333 16175 26367
rect 16117 26327 16175 26333
rect 18690 26324 18696 26376
rect 18748 26324 18754 26376
rect 19978 26324 19984 26376
rect 20036 26324 20042 26376
rect 20438 26324 20444 26376
rect 20496 26324 20502 26376
rect 22066 26364 22094 26540
rect 24412 26441 24440 26540
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 25774 26460 25780 26512
rect 25832 26460 25838 26512
rect 24397 26435 24455 26441
rect 24397 26401 24409 26435
rect 24443 26401 24455 26435
rect 24397 26395 24455 26401
rect 20640 26336 22094 26364
rect 16025 26299 16083 26305
rect 16025 26296 16037 26299
rect 15304 26268 16037 26296
rect 14093 26259 14151 26265
rect 16025 26265 16037 26268
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 17865 26299 17923 26305
rect 17865 26265 17877 26299
rect 17911 26265 17923 26299
rect 19996 26296 20024 26324
rect 20640 26296 20668 26336
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 19996 26268 20668 26296
rect 20708 26299 20766 26305
rect 17865 26259 17923 26265
rect 20708 26265 20720 26299
rect 20754 26296 20766 26299
rect 21358 26296 21364 26308
rect 20754 26268 21364 26296
rect 20754 26265 20766 26268
rect 20708 26259 20766 26265
rect 8757 26231 8815 26237
rect 8757 26197 8769 26231
rect 8803 26197 8815 26231
rect 8757 26191 8815 26197
rect 10410 26188 10416 26240
rect 10468 26188 10474 26240
rect 11698 26188 11704 26240
rect 11756 26188 11762 26240
rect 12894 26188 12900 26240
rect 12952 26228 12958 26240
rect 13081 26231 13139 26237
rect 13081 26228 13093 26231
rect 12952 26200 13093 26228
rect 12952 26188 12958 26200
rect 13081 26197 13093 26200
rect 13127 26197 13139 26231
rect 17880 26228 17908 26259
rect 21358 26256 21364 26268
rect 21416 26256 21422 26308
rect 24642 26299 24700 26305
rect 24642 26296 24654 26299
rect 24228 26268 24654 26296
rect 17954 26228 17960 26240
rect 17880 26200 17960 26228
rect 13081 26191 13139 26197
rect 17954 26188 17960 26200
rect 18012 26188 18018 26240
rect 24228 26237 24256 26268
rect 24642 26265 24654 26268
rect 24688 26265 24700 26299
rect 24642 26259 24700 26265
rect 24213 26231 24271 26237
rect 24213 26197 24225 26231
rect 24259 26197 24271 26231
rect 24213 26191 24271 26197
rect 1104 26138 31280 26160
rect 1104 26086 4922 26138
rect 4974 26086 4986 26138
rect 5038 26086 5050 26138
rect 5102 26086 5114 26138
rect 5166 26086 5178 26138
rect 5230 26086 5242 26138
rect 5294 26086 10922 26138
rect 10974 26086 10986 26138
rect 11038 26086 11050 26138
rect 11102 26086 11114 26138
rect 11166 26086 11178 26138
rect 11230 26086 11242 26138
rect 11294 26086 16922 26138
rect 16974 26086 16986 26138
rect 17038 26086 17050 26138
rect 17102 26086 17114 26138
rect 17166 26086 17178 26138
rect 17230 26086 17242 26138
rect 17294 26086 22922 26138
rect 22974 26086 22986 26138
rect 23038 26086 23050 26138
rect 23102 26086 23114 26138
rect 23166 26086 23178 26138
rect 23230 26086 23242 26138
rect 23294 26086 28922 26138
rect 28974 26086 28986 26138
rect 29038 26086 29050 26138
rect 29102 26086 29114 26138
rect 29166 26086 29178 26138
rect 29230 26086 29242 26138
rect 29294 26086 31280 26138
rect 1104 26064 31280 26086
rect 8570 25984 8576 26036
rect 8628 26024 8634 26036
rect 9309 26027 9367 26033
rect 9309 26024 9321 26027
rect 8628 25996 9321 26024
rect 8628 25984 8634 25996
rect 9309 25993 9321 25996
rect 9355 25993 9367 26027
rect 9309 25987 9367 25993
rect 9677 26027 9735 26033
rect 9677 25993 9689 26027
rect 9723 26024 9735 26027
rect 10042 26024 10048 26036
rect 9723 25996 10048 26024
rect 9723 25993 9735 25996
rect 9677 25987 9735 25993
rect 10042 25984 10048 25996
rect 10100 25984 10106 26036
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10505 26027 10563 26033
rect 10505 26024 10517 26027
rect 10468 25996 10517 26024
rect 10468 25984 10474 25996
rect 10505 25993 10517 25996
rect 10551 25993 10563 26027
rect 10505 25987 10563 25993
rect 12805 26027 12863 26033
rect 12805 25993 12817 26027
rect 12851 26024 12863 26027
rect 14277 26027 14335 26033
rect 12851 25996 13032 26024
rect 12851 25993 12863 25996
rect 12805 25987 12863 25993
rect 10597 25959 10655 25965
rect 10597 25956 10609 25959
rect 9692 25928 10609 25956
rect 9692 25900 9720 25928
rect 10597 25925 10609 25928
rect 10643 25925 10655 25959
rect 10597 25919 10655 25925
rect 12894 25916 12900 25968
rect 12952 25916 12958 25968
rect 13004 25956 13032 25996
rect 14277 25993 14289 26027
rect 14323 26024 14335 26027
rect 14642 26024 14648 26036
rect 14323 25996 14648 26024
rect 14323 25993 14335 25996
rect 14277 25987 14335 25993
rect 14642 25984 14648 25996
rect 14700 25984 14706 26036
rect 24026 25984 24032 26036
rect 24084 26024 24090 26036
rect 24213 26027 24271 26033
rect 24213 26024 24225 26027
rect 24084 25996 24225 26024
rect 24084 25984 24090 25996
rect 24213 25993 24225 25996
rect 24259 25993 24271 26027
rect 24213 25987 24271 25993
rect 13164 25959 13222 25965
rect 13164 25956 13176 25959
rect 13004 25928 13176 25956
rect 13164 25925 13176 25928
rect 13210 25925 13222 25959
rect 13164 25919 13222 25925
rect 19978 25916 19984 25968
rect 20036 25916 20042 25968
rect 7374 25848 7380 25900
rect 7432 25888 7438 25900
rect 8110 25897 8116 25900
rect 7837 25891 7895 25897
rect 7837 25888 7849 25891
rect 7432 25860 7849 25888
rect 7432 25848 7438 25860
rect 7837 25857 7849 25860
rect 7883 25857 7895 25891
rect 7837 25851 7895 25857
rect 8104 25851 8116 25897
rect 8110 25848 8116 25851
rect 8168 25848 8174 25900
rect 9674 25848 9680 25900
rect 9732 25848 9738 25900
rect 9769 25891 9827 25897
rect 9769 25857 9781 25891
rect 9815 25888 9827 25891
rect 12434 25888 12440 25900
rect 9815 25860 12440 25888
rect 9815 25857 9827 25860
rect 9769 25851 9827 25857
rect 5534 25780 5540 25832
rect 5592 25780 5598 25832
rect 9784 25820 9812 25851
rect 12434 25848 12440 25860
rect 12492 25848 12498 25900
rect 12621 25891 12679 25897
rect 12621 25857 12633 25891
rect 12667 25888 12679 25891
rect 12912 25888 12940 25916
rect 12667 25860 12940 25888
rect 12667 25857 12679 25860
rect 12621 25851 12679 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 19153 25891 19211 25897
rect 19153 25888 19165 25891
rect 18012 25860 19165 25888
rect 18012 25848 18018 25860
rect 19153 25857 19165 25860
rect 19199 25857 19211 25891
rect 19153 25851 19211 25857
rect 24581 25891 24639 25897
rect 24581 25857 24593 25891
rect 24627 25888 24639 25891
rect 25041 25891 25099 25897
rect 25041 25888 25053 25891
rect 24627 25860 25053 25888
rect 24627 25857 24639 25860
rect 24581 25851 24639 25857
rect 25041 25857 25053 25860
rect 25087 25857 25099 25891
rect 25041 25851 25099 25857
rect 25685 25891 25743 25897
rect 25685 25857 25697 25891
rect 25731 25888 25743 25891
rect 25774 25888 25780 25900
rect 25731 25860 25780 25888
rect 25731 25857 25743 25860
rect 25685 25851 25743 25857
rect 25774 25848 25780 25860
rect 25832 25848 25838 25900
rect 8864 25792 9812 25820
rect 8864 25696 8892 25792
rect 9950 25780 9956 25832
rect 10008 25780 10014 25832
rect 10594 25780 10600 25832
rect 10652 25820 10658 25832
rect 10689 25823 10747 25829
rect 10689 25820 10701 25823
rect 10652 25792 10701 25820
rect 10652 25780 10658 25792
rect 10689 25789 10701 25792
rect 10735 25789 10747 25823
rect 10689 25783 10747 25789
rect 12342 25780 12348 25832
rect 12400 25820 12406 25832
rect 12526 25820 12532 25832
rect 12400 25792 12532 25820
rect 12400 25780 12406 25792
rect 12526 25780 12532 25792
rect 12584 25820 12590 25832
rect 12897 25823 12955 25829
rect 12897 25820 12909 25823
rect 12584 25792 12909 25820
rect 12584 25780 12590 25792
rect 12897 25789 12909 25792
rect 12943 25789 12955 25823
rect 12897 25783 12955 25789
rect 20254 25780 20260 25832
rect 20312 25780 20318 25832
rect 24486 25780 24492 25832
rect 24544 25820 24550 25832
rect 24673 25823 24731 25829
rect 24673 25820 24685 25823
rect 24544 25792 24685 25820
rect 24544 25780 24550 25792
rect 24673 25789 24685 25792
rect 24719 25789 24731 25823
rect 24673 25783 24731 25789
rect 24765 25823 24823 25829
rect 24765 25789 24777 25823
rect 24811 25820 24823 25823
rect 24854 25820 24860 25832
rect 24811 25792 24860 25820
rect 24811 25789 24823 25792
rect 24765 25783 24823 25789
rect 9217 25755 9275 25761
rect 9217 25721 9229 25755
rect 9263 25752 9275 25755
rect 10502 25752 10508 25764
rect 9263 25724 10508 25752
rect 9263 25721 9275 25724
rect 9217 25715 9275 25721
rect 10502 25712 10508 25724
rect 10560 25712 10566 25764
rect 20272 25752 20300 25780
rect 24780 25752 24808 25783
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 20272 25724 24808 25752
rect 4890 25644 4896 25696
rect 4948 25644 4954 25696
rect 7006 25644 7012 25696
rect 7064 25684 7070 25696
rect 8846 25684 8852 25696
rect 7064 25656 8852 25684
rect 7064 25644 7070 25656
rect 8846 25644 8852 25656
rect 8904 25644 8910 25696
rect 9306 25644 9312 25696
rect 9364 25684 9370 25696
rect 10137 25687 10195 25693
rect 10137 25684 10149 25687
rect 9364 25656 10149 25684
rect 9364 25644 9370 25656
rect 10137 25653 10149 25656
rect 10183 25653 10195 25687
rect 10137 25647 10195 25653
rect 11974 25644 11980 25696
rect 12032 25684 12038 25696
rect 13078 25684 13084 25696
rect 12032 25656 13084 25684
rect 12032 25644 12038 25656
rect 13078 25644 13084 25656
rect 13136 25684 13142 25696
rect 14734 25684 14740 25696
rect 13136 25656 14740 25684
rect 13136 25644 13142 25656
rect 14734 25644 14740 25656
rect 14792 25644 14798 25696
rect 1104 25594 31280 25616
rect 1104 25542 4182 25594
rect 4234 25542 4246 25594
rect 4298 25542 4310 25594
rect 4362 25542 4374 25594
rect 4426 25542 4438 25594
rect 4490 25542 4502 25594
rect 4554 25542 10182 25594
rect 10234 25542 10246 25594
rect 10298 25542 10310 25594
rect 10362 25542 10374 25594
rect 10426 25542 10438 25594
rect 10490 25542 10502 25594
rect 10554 25542 16182 25594
rect 16234 25542 16246 25594
rect 16298 25542 16310 25594
rect 16362 25542 16374 25594
rect 16426 25542 16438 25594
rect 16490 25542 16502 25594
rect 16554 25542 22182 25594
rect 22234 25542 22246 25594
rect 22298 25542 22310 25594
rect 22362 25542 22374 25594
rect 22426 25542 22438 25594
rect 22490 25542 22502 25594
rect 22554 25542 28182 25594
rect 28234 25542 28246 25594
rect 28298 25542 28310 25594
rect 28362 25542 28374 25594
rect 28426 25542 28438 25594
rect 28490 25542 28502 25594
rect 28554 25542 31280 25594
rect 1104 25520 31280 25542
rect 4890 25480 4896 25492
rect 4632 25452 4896 25480
rect 4632 25285 4660 25452
rect 4890 25440 4896 25452
rect 4948 25440 4954 25492
rect 5350 25480 5356 25492
rect 5092 25452 5356 25480
rect 4893 25347 4951 25353
rect 4893 25313 4905 25347
rect 4939 25344 4951 25347
rect 5092 25344 5120 25452
rect 5350 25440 5356 25452
rect 5408 25480 5414 25492
rect 5994 25480 6000 25492
rect 5408 25452 6000 25480
rect 5408 25440 5414 25452
rect 5994 25440 6000 25452
rect 6052 25440 6058 25492
rect 7374 25480 7380 25492
rect 6288 25452 7380 25480
rect 4939 25316 5120 25344
rect 4939 25313 4951 25316
rect 4893 25307 4951 25313
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25276 4215 25279
rect 4617 25279 4675 25285
rect 4203 25248 4292 25276
rect 4203 25245 4215 25248
rect 4157 25239 4215 25245
rect 3970 25100 3976 25152
rect 4028 25100 4034 25152
rect 4264 25149 4292 25248
rect 4617 25245 4629 25279
rect 4663 25245 4675 25279
rect 4617 25239 4675 25245
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 5077 25279 5135 25285
rect 5077 25276 5089 25279
rect 4764 25248 5089 25276
rect 4764 25236 4770 25248
rect 5077 25245 5089 25248
rect 5123 25276 5135 25279
rect 6288 25276 6316 25452
rect 7374 25440 7380 25452
rect 7432 25440 7438 25492
rect 8110 25440 8116 25492
rect 8168 25480 8174 25492
rect 8205 25483 8263 25489
rect 8205 25480 8217 25483
rect 8168 25452 8217 25480
rect 8168 25440 8174 25452
rect 8205 25449 8217 25452
rect 8251 25449 8263 25483
rect 8205 25443 8263 25449
rect 9306 25440 9312 25492
rect 9364 25440 9370 25492
rect 9582 25440 9588 25492
rect 9640 25480 9646 25492
rect 12342 25480 12348 25492
rect 9640 25452 12348 25480
rect 9640 25440 9646 25452
rect 12342 25440 12348 25452
rect 12400 25440 12406 25492
rect 30837 25483 30895 25489
rect 30837 25449 30849 25483
rect 30883 25480 30895 25483
rect 30883 25452 31340 25480
rect 30883 25449 30895 25452
rect 30837 25443 30895 25449
rect 6457 25415 6515 25421
rect 6457 25381 6469 25415
rect 6503 25412 6515 25415
rect 6638 25412 6644 25424
rect 6503 25384 6644 25412
rect 6503 25381 6515 25384
rect 6457 25375 6515 25381
rect 6638 25372 6644 25384
rect 6696 25412 6702 25424
rect 6696 25384 7972 25412
rect 6696 25372 6702 25384
rect 7193 25347 7251 25353
rect 7193 25313 7205 25347
rect 7239 25344 7251 25347
rect 7466 25344 7472 25356
rect 7239 25316 7472 25344
rect 7239 25313 7251 25316
rect 7193 25307 7251 25313
rect 5123 25248 6316 25276
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 5344 25211 5402 25217
rect 5344 25177 5356 25211
rect 5390 25208 5402 25211
rect 5442 25208 5448 25220
rect 5390 25180 5448 25208
rect 5390 25177 5402 25180
rect 5344 25171 5402 25177
rect 5442 25168 5448 25180
rect 5500 25168 5506 25220
rect 6822 25168 6828 25220
rect 6880 25208 6886 25220
rect 7208 25208 7236 25307
rect 7466 25304 7472 25316
rect 7524 25304 7530 25356
rect 7944 25353 7972 25384
rect 7929 25347 7987 25353
rect 7929 25313 7941 25347
rect 7975 25313 7987 25347
rect 9324 25344 9352 25440
rect 9600 25353 9628 25440
rect 31312 25424 31340 25452
rect 10965 25415 11023 25421
rect 10965 25381 10977 25415
rect 11011 25412 11023 25415
rect 11011 25384 11652 25412
rect 11011 25381 11023 25384
rect 10965 25375 11023 25381
rect 11624 25356 11652 25384
rect 31294 25372 31300 25424
rect 31352 25372 31358 25424
rect 7929 25307 7987 25313
rect 8404 25316 9352 25344
rect 9585 25347 9643 25353
rect 8404 25285 8432 25316
rect 9585 25313 9597 25347
rect 9631 25313 9643 25347
rect 9585 25307 9643 25313
rect 11606 25304 11612 25356
rect 11664 25304 11670 25356
rect 17862 25304 17868 25356
rect 17920 25344 17926 25356
rect 18049 25347 18107 25353
rect 18049 25344 18061 25347
rect 17920 25316 18061 25344
rect 17920 25304 17926 25316
rect 18049 25313 18061 25316
rect 18095 25313 18107 25347
rect 18049 25307 18107 25313
rect 18874 25304 18880 25356
rect 18932 25304 18938 25356
rect 8389 25279 8447 25285
rect 8389 25245 8401 25279
rect 8435 25245 8447 25279
rect 8389 25239 8447 25245
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25276 12127 25279
rect 14737 25279 14795 25285
rect 12115 25248 12572 25276
rect 12115 25245 12127 25248
rect 12069 25239 12127 25245
rect 12342 25217 12348 25220
rect 9830 25211 9888 25217
rect 9830 25208 9842 25211
rect 6880 25180 7236 25208
rect 9508 25180 9842 25208
rect 6880 25168 6886 25180
rect 4249 25143 4307 25149
rect 4249 25109 4261 25143
rect 4295 25109 4307 25143
rect 4249 25103 4307 25109
rect 4709 25143 4767 25149
rect 4709 25109 4721 25143
rect 4755 25140 4767 25143
rect 4798 25140 4804 25152
rect 4755 25112 4804 25140
rect 4755 25109 4767 25112
rect 4709 25103 4767 25109
rect 4798 25100 4804 25112
rect 4856 25100 4862 25152
rect 6086 25100 6092 25152
rect 6144 25140 6150 25152
rect 6549 25143 6607 25149
rect 6549 25140 6561 25143
rect 6144 25112 6561 25140
rect 6144 25100 6150 25112
rect 6549 25109 6561 25112
rect 6595 25109 6607 25143
rect 6549 25103 6607 25109
rect 6914 25100 6920 25152
rect 6972 25100 6978 25152
rect 9508 25149 9536 25180
rect 9830 25177 9842 25180
rect 9876 25177 9888 25211
rect 9830 25171 9888 25177
rect 12336 25171 12348 25217
rect 12342 25168 12348 25171
rect 12400 25168 12406 25220
rect 12544 25152 12572 25248
rect 14737 25245 14749 25279
rect 14783 25245 14795 25279
rect 14737 25239 14795 25245
rect 17957 25279 18015 25285
rect 17957 25245 17969 25279
rect 18003 25276 18015 25279
rect 18003 25248 19748 25276
rect 18003 25245 18015 25248
rect 17957 25239 18015 25245
rect 14752 25208 14780 25239
rect 13464 25180 14780 25208
rect 17865 25211 17923 25217
rect 13464 25152 13492 25180
rect 17865 25177 17877 25211
rect 17911 25208 17923 25211
rect 18414 25208 18420 25220
rect 17911 25180 18420 25208
rect 17911 25177 17923 25180
rect 17865 25171 17923 25177
rect 18414 25168 18420 25180
rect 18472 25168 18478 25220
rect 18693 25211 18751 25217
rect 18693 25177 18705 25211
rect 18739 25208 18751 25211
rect 19245 25211 19303 25217
rect 19245 25208 19257 25211
rect 18739 25180 19257 25208
rect 18739 25177 18751 25180
rect 18693 25171 18751 25177
rect 19245 25177 19257 25180
rect 19291 25177 19303 25211
rect 19720 25208 19748 25248
rect 19794 25236 19800 25288
rect 19852 25236 19858 25288
rect 30650 25236 30656 25288
rect 30708 25236 30714 25288
rect 20806 25208 20812 25220
rect 19720 25180 20812 25208
rect 19245 25171 19303 25177
rect 20806 25168 20812 25180
rect 20864 25168 20870 25220
rect 7009 25143 7067 25149
rect 7009 25109 7021 25143
rect 7055 25140 7067 25143
rect 7377 25143 7435 25149
rect 7377 25140 7389 25143
rect 7055 25112 7389 25140
rect 7055 25109 7067 25112
rect 7009 25103 7067 25109
rect 7377 25109 7389 25112
rect 7423 25109 7435 25143
rect 7377 25103 7435 25109
rect 9493 25143 9551 25149
rect 9493 25109 9505 25143
rect 9539 25109 9551 25143
rect 9493 25103 9551 25109
rect 9950 25100 9956 25152
rect 10008 25140 10014 25152
rect 11057 25143 11115 25149
rect 11057 25140 11069 25143
rect 10008 25112 11069 25140
rect 10008 25100 10014 25112
rect 11057 25109 11069 25112
rect 11103 25109 11115 25143
rect 11057 25103 11115 25109
rect 12526 25100 12532 25152
rect 12584 25100 12590 25152
rect 13446 25100 13452 25152
rect 13504 25100 13510 25152
rect 14090 25100 14096 25152
rect 14148 25100 14154 25152
rect 17494 25100 17500 25152
rect 17552 25100 17558 25152
rect 18322 25100 18328 25152
rect 18380 25100 18386 25152
rect 18785 25143 18843 25149
rect 18785 25109 18797 25143
rect 18831 25140 18843 25143
rect 20622 25140 20628 25152
rect 18831 25112 20628 25140
rect 18831 25109 18843 25112
rect 18785 25103 18843 25109
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 1104 25050 31280 25072
rect 1104 24998 4922 25050
rect 4974 24998 4986 25050
rect 5038 24998 5050 25050
rect 5102 24998 5114 25050
rect 5166 24998 5178 25050
rect 5230 24998 5242 25050
rect 5294 24998 10922 25050
rect 10974 24998 10986 25050
rect 11038 24998 11050 25050
rect 11102 24998 11114 25050
rect 11166 24998 11178 25050
rect 11230 24998 11242 25050
rect 11294 24998 16922 25050
rect 16974 24998 16986 25050
rect 17038 24998 17050 25050
rect 17102 24998 17114 25050
rect 17166 24998 17178 25050
rect 17230 24998 17242 25050
rect 17294 24998 22922 25050
rect 22974 24998 22986 25050
rect 23038 24998 23050 25050
rect 23102 24998 23114 25050
rect 23166 24998 23178 25050
rect 23230 24998 23242 25050
rect 23294 24998 28922 25050
rect 28974 24998 28986 25050
rect 29038 24998 29050 25050
rect 29102 24998 29114 25050
rect 29166 24998 29178 25050
rect 29230 24998 29242 25050
rect 29294 24998 31280 25050
rect 1104 24976 31280 24998
rect 4706 24936 4712 24948
rect 3896 24908 4712 24936
rect 3697 24803 3755 24809
rect 3697 24769 3709 24803
rect 3743 24800 3755 24803
rect 3896 24800 3924 24908
rect 4706 24896 4712 24908
rect 4764 24896 4770 24948
rect 5442 24896 5448 24948
rect 5500 24896 5506 24948
rect 5552 24908 8248 24936
rect 4798 24828 4804 24880
rect 4856 24868 4862 24880
rect 5552 24868 5580 24908
rect 6086 24868 6092 24880
rect 4856 24840 5580 24868
rect 5644 24840 6092 24868
rect 4856 24828 4862 24840
rect 3970 24809 3976 24812
rect 3743 24772 3924 24800
rect 3743 24769 3755 24772
rect 3697 24763 3755 24769
rect 3964 24763 3976 24809
rect 4028 24800 4034 24812
rect 5644 24809 5672 24840
rect 6086 24828 6092 24840
rect 6144 24828 6150 24880
rect 6638 24828 6644 24880
rect 6696 24828 6702 24880
rect 7374 24828 7380 24880
rect 7432 24868 7438 24880
rect 8110 24868 8116 24880
rect 7432 24840 8116 24868
rect 7432 24828 7438 24840
rect 8110 24828 8116 24840
rect 8168 24828 8174 24880
rect 8220 24868 8248 24908
rect 9306 24896 9312 24948
rect 9364 24936 9370 24948
rect 9585 24939 9643 24945
rect 9585 24936 9597 24939
rect 9364 24908 9597 24936
rect 9364 24896 9370 24908
rect 9585 24905 9597 24908
rect 9631 24905 9643 24939
rect 9585 24899 9643 24905
rect 9950 24896 9956 24948
rect 10008 24896 10014 24948
rect 12253 24939 12311 24945
rect 12253 24905 12265 24939
rect 12299 24936 12311 24939
rect 12342 24936 12348 24948
rect 12299 24908 12348 24936
rect 12299 24905 12311 24908
rect 12253 24899 12311 24905
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 12434 24896 12440 24948
rect 12492 24936 12498 24948
rect 12897 24939 12955 24945
rect 12492 24908 12848 24936
rect 12492 24896 12498 24908
rect 9674 24868 9680 24880
rect 8220 24840 9680 24868
rect 9674 24828 9680 24840
rect 9732 24828 9738 24880
rect 11241 24871 11299 24877
rect 11241 24837 11253 24871
rect 11287 24868 11299 24871
rect 12526 24868 12532 24880
rect 11287 24840 12532 24868
rect 11287 24837 11299 24840
rect 11241 24831 11299 24837
rect 12526 24828 12532 24840
rect 12584 24828 12590 24880
rect 5629 24803 5687 24809
rect 4028 24772 4064 24800
rect 3970 24760 3976 24763
rect 4028 24760 4034 24772
rect 5629 24769 5641 24803
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 6365 24803 6423 24809
rect 6365 24769 6377 24803
rect 6411 24769 6423 24803
rect 6365 24763 6423 24769
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 6733 24803 6791 24809
rect 6733 24769 6745 24803
rect 6779 24800 6791 24803
rect 7650 24800 7656 24812
rect 6779 24772 7656 24800
rect 6779 24769 6791 24772
rect 6733 24763 6791 24769
rect 5077 24667 5135 24673
rect 5077 24633 5089 24667
rect 5123 24664 5135 24667
rect 5534 24664 5540 24676
rect 5123 24636 5540 24664
rect 5123 24633 5135 24636
rect 5077 24627 5135 24633
rect 5534 24624 5540 24636
rect 5592 24664 5598 24676
rect 6380 24664 6408 24763
rect 6564 24732 6592 24763
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 8941 24803 8999 24809
rect 8941 24769 8953 24803
rect 8987 24800 8999 24803
rect 10413 24803 10471 24809
rect 10413 24800 10425 24803
rect 8987 24772 10425 24800
rect 8987 24769 8999 24772
rect 8941 24763 8999 24769
rect 10413 24769 10425 24772
rect 10459 24800 10471 24803
rect 10686 24800 10692 24812
rect 10459 24772 10692 24800
rect 10459 24769 10471 24772
rect 10413 24763 10471 24769
rect 10686 24760 10692 24772
rect 10744 24760 10750 24812
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24800 11575 24803
rect 11606 24800 11612 24812
rect 11563 24772 11612 24800
rect 11563 24769 11575 24772
rect 11517 24763 11575 24769
rect 11606 24760 11612 24772
rect 11664 24760 11670 24812
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 11793 24803 11851 24809
rect 11793 24769 11805 24803
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 12158 24800 12164 24812
rect 11931 24772 12164 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 7190 24732 7196 24744
rect 6564 24704 7196 24732
rect 7190 24692 7196 24704
rect 7248 24692 7254 24744
rect 9674 24692 9680 24744
rect 9732 24732 9738 24744
rect 10045 24735 10103 24741
rect 10045 24732 10057 24735
rect 9732 24704 10057 24732
rect 9732 24692 9738 24704
rect 10045 24701 10057 24704
rect 10091 24701 10103 24735
rect 10045 24695 10103 24701
rect 10134 24692 10140 24744
rect 10192 24692 10198 24744
rect 5592 24636 6408 24664
rect 5592 24624 5598 24636
rect 6914 24556 6920 24608
rect 6972 24556 6978 24608
rect 11422 24556 11428 24608
rect 11480 24596 11486 24608
rect 11716 24596 11744 24763
rect 11808 24664 11836 24763
rect 12158 24760 12164 24772
rect 12216 24760 12222 24812
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24800 12495 24803
rect 12820 24800 12848 24908
rect 12897 24905 12909 24939
rect 12943 24936 12955 24939
rect 14090 24936 14096 24948
rect 12943 24908 14096 24936
rect 12943 24905 12955 24908
rect 12897 24899 12955 24905
rect 14090 24896 14096 24908
rect 14148 24896 14154 24948
rect 14642 24896 14648 24948
rect 14700 24896 14706 24948
rect 17494 24896 17500 24948
rect 17552 24896 17558 24948
rect 18414 24896 18420 24948
rect 18472 24936 18478 24948
rect 18969 24939 19027 24945
rect 18969 24936 18981 24939
rect 18472 24908 18981 24936
rect 18472 24896 18478 24908
rect 18969 24905 18981 24908
rect 19015 24905 19027 24939
rect 18969 24899 19027 24905
rect 14660 24868 14688 24896
rect 13740 24840 14688 24868
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12483 24772 12572 24800
rect 12820 24772 13001 24800
rect 12483 24769 12495 24772
rect 12437 24763 12495 24769
rect 12544 24673 12572 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13538 24760 13544 24812
rect 13596 24760 13602 24812
rect 13740 24809 13768 24840
rect 13725 24803 13783 24809
rect 13725 24769 13737 24803
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 13817 24803 13875 24809
rect 13817 24769 13829 24803
rect 13863 24769 13875 24803
rect 13817 24763 13875 24769
rect 17405 24803 17463 24809
rect 17405 24769 17417 24803
rect 17451 24800 17463 24803
rect 17512 24800 17540 24896
rect 19610 24828 19616 24880
rect 19668 24868 19674 24880
rect 20717 24871 20775 24877
rect 19668 24840 19840 24868
rect 19668 24828 19674 24840
rect 17451 24772 17540 24800
rect 17451 24769 17463 24772
rect 17405 24763 17463 24769
rect 13173 24735 13231 24741
rect 13173 24701 13185 24735
rect 13219 24732 13231 24735
rect 13832 24732 13860 24763
rect 17586 24760 17592 24812
rect 17644 24800 17650 24812
rect 17753 24803 17811 24809
rect 17753 24800 17765 24803
rect 17644 24772 17765 24800
rect 17644 24760 17650 24772
rect 17753 24769 17765 24772
rect 17799 24769 17811 24803
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 17753 24763 17811 24769
rect 19536 24772 19717 24800
rect 13219 24704 13676 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 12529 24667 12587 24673
rect 11808 24636 12434 24664
rect 11974 24596 11980 24608
rect 11480 24568 11980 24596
rect 11480 24556 11486 24568
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12066 24556 12072 24608
rect 12124 24556 12130 24608
rect 12406 24596 12434 24636
rect 12529 24633 12541 24667
rect 12575 24633 12587 24667
rect 13446 24664 13452 24676
rect 12529 24627 12587 24633
rect 12636 24636 13452 24664
rect 12636 24596 12664 24636
rect 13446 24624 13452 24636
rect 13504 24624 13510 24676
rect 12406 24568 12664 24596
rect 13354 24556 13360 24608
rect 13412 24556 13418 24608
rect 13648 24596 13676 24704
rect 13740 24704 13860 24732
rect 13740 24676 13768 24704
rect 14550 24692 14556 24744
rect 14608 24692 14614 24744
rect 14918 24692 14924 24744
rect 14976 24692 14982 24744
rect 19536 24741 19564 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19812 24800 19840 24840
rect 20717 24837 20729 24871
rect 20763 24868 20775 24871
rect 21821 24871 21879 24877
rect 21821 24868 21833 24871
rect 20763 24840 21833 24868
rect 20763 24837 20775 24840
rect 20717 24831 20775 24837
rect 21821 24837 21833 24840
rect 21867 24837 21879 24871
rect 21821 24831 21879 24837
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 19812 24772 19901 24800
rect 19705 24763 19763 24769
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 19981 24803 20039 24809
rect 19981 24769 19993 24803
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24800 20131 24803
rect 20346 24800 20352 24812
rect 20119 24772 20352 24800
rect 20119 24769 20131 24772
rect 20073 24763 20131 24769
rect 17497 24735 17555 24741
rect 17497 24701 17509 24735
rect 17543 24701 17555 24735
rect 17497 24695 17555 24701
rect 19521 24735 19579 24741
rect 19521 24701 19533 24735
rect 19567 24701 19579 24735
rect 19521 24695 19579 24701
rect 13722 24624 13728 24676
rect 13780 24624 13786 24676
rect 14568 24664 14596 24692
rect 13832 24636 14596 24664
rect 13832 24596 13860 24636
rect 17512 24608 17540 24695
rect 19536 24664 19564 24695
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 19996 24732 20024 24763
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20806 24760 20812 24812
rect 20864 24760 20870 24812
rect 21358 24760 21364 24812
rect 21416 24760 21422 24812
rect 19852 24704 20024 24732
rect 19852 24692 19858 24704
rect 18432 24636 19564 24664
rect 18432 24608 18460 24636
rect 13648 24568 13860 24596
rect 14366 24556 14372 24608
rect 14424 24556 14430 24608
rect 17218 24556 17224 24608
rect 17276 24556 17282 24608
rect 17494 24556 17500 24608
rect 17552 24556 17558 24608
rect 18414 24556 18420 24608
rect 18472 24556 18478 24608
rect 18877 24599 18935 24605
rect 18877 24565 18889 24599
rect 18923 24596 18935 24599
rect 19812 24596 19840 24692
rect 19886 24624 19892 24676
rect 19944 24664 19950 24676
rect 20349 24667 20407 24673
rect 20349 24664 20361 24667
rect 19944 24636 20361 24664
rect 19944 24624 19950 24636
rect 20349 24633 20361 24636
rect 20395 24633 20407 24667
rect 20824 24664 20852 24760
rect 20898 24692 20904 24744
rect 20956 24692 20962 24744
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 21324 24704 22385 24732
rect 21324 24692 21330 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 24394 24692 24400 24744
rect 24452 24692 24458 24744
rect 25222 24692 25228 24744
rect 25280 24692 25286 24744
rect 23566 24664 23572 24676
rect 20824 24636 23572 24664
rect 20349 24627 20407 24633
rect 23566 24624 23572 24636
rect 23624 24624 23630 24676
rect 24670 24664 24676 24676
rect 23768 24636 24676 24664
rect 18923 24568 19840 24596
rect 18923 24565 18935 24568
rect 18877 24559 18935 24565
rect 20254 24556 20260 24608
rect 20312 24556 20318 24608
rect 21174 24556 21180 24608
rect 21232 24556 21238 24608
rect 22094 24556 22100 24608
rect 22152 24596 22158 24608
rect 23768 24596 23796 24636
rect 24670 24624 24676 24636
rect 24728 24624 24734 24676
rect 22152 24568 23796 24596
rect 22152 24556 22158 24568
rect 23842 24556 23848 24608
rect 23900 24556 23906 24608
rect 24578 24556 24584 24608
rect 24636 24556 24642 24608
rect 1104 24506 31280 24528
rect 1104 24454 4182 24506
rect 4234 24454 4246 24506
rect 4298 24454 4310 24506
rect 4362 24454 4374 24506
rect 4426 24454 4438 24506
rect 4490 24454 4502 24506
rect 4554 24454 10182 24506
rect 10234 24454 10246 24506
rect 10298 24454 10310 24506
rect 10362 24454 10374 24506
rect 10426 24454 10438 24506
rect 10490 24454 10502 24506
rect 10554 24454 16182 24506
rect 16234 24454 16246 24506
rect 16298 24454 16310 24506
rect 16362 24454 16374 24506
rect 16426 24454 16438 24506
rect 16490 24454 16502 24506
rect 16554 24454 22182 24506
rect 22234 24454 22246 24506
rect 22298 24454 22310 24506
rect 22362 24454 22374 24506
rect 22426 24454 22438 24506
rect 22490 24454 22502 24506
rect 22554 24454 28182 24506
rect 28234 24454 28246 24506
rect 28298 24454 28310 24506
rect 28362 24454 28374 24506
rect 28426 24454 28438 24506
rect 28490 24454 28502 24506
rect 28554 24454 31280 24506
rect 1104 24432 31280 24454
rect 6914 24352 6920 24404
rect 6972 24352 6978 24404
rect 11977 24395 12035 24401
rect 11977 24361 11989 24395
rect 12023 24392 12035 24395
rect 12066 24392 12072 24404
rect 12023 24364 12072 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 13354 24392 13360 24404
rect 12406 24364 13360 24392
rect 6932 24256 6960 24352
rect 11885 24259 11943 24265
rect 6932 24228 11836 24256
rect 8570 24148 8576 24200
rect 8628 24148 8634 24200
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24188 10379 24191
rect 10778 24188 10784 24200
rect 10367 24160 10784 24188
rect 10367 24157 10379 24160
rect 10321 24151 10379 24157
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 11698 24148 11704 24200
rect 11756 24148 11762 24200
rect 11808 24188 11836 24228
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 12406 24256 12434 24364
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 14918 24392 14924 24404
rect 14323 24364 14924 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 18414 24352 18420 24404
rect 18472 24352 18478 24404
rect 19886 24352 19892 24404
rect 19944 24352 19950 24404
rect 20162 24352 20168 24404
rect 20220 24392 20226 24404
rect 20220 24364 20852 24392
rect 20220 24352 20226 24364
rect 11931 24228 12434 24256
rect 15657 24259 15715 24265
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 15657 24225 15669 24259
rect 15703 24256 15715 24259
rect 16114 24256 16120 24268
rect 15703 24228 16120 24256
rect 15703 24225 15715 24228
rect 15657 24219 15715 24225
rect 16114 24216 16120 24228
rect 16172 24256 16178 24268
rect 19904 24256 19932 24352
rect 20824 24324 20852 24364
rect 21266 24352 21272 24404
rect 21324 24352 21330 24404
rect 21358 24352 21364 24404
rect 21416 24352 21422 24404
rect 24029 24395 24087 24401
rect 22572 24364 23612 24392
rect 22094 24324 22100 24336
rect 20824 24296 22100 24324
rect 22094 24284 22100 24296
rect 22152 24284 22158 24336
rect 16172 24228 17080 24256
rect 16172 24216 16178 24228
rect 11977 24191 12035 24197
rect 11977 24188 11989 24191
rect 11808 24160 11989 24188
rect 11977 24157 11989 24160
rect 12023 24157 12035 24191
rect 11977 24151 12035 24157
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 17052 24197 17080 24228
rect 19628 24228 19932 24256
rect 19628 24197 19656 24228
rect 20990 24216 20996 24268
rect 21048 24256 21054 24268
rect 21913 24259 21971 24265
rect 21913 24256 21925 24259
rect 21048 24228 21925 24256
rect 21048 24216 21054 24228
rect 21913 24225 21925 24228
rect 21959 24225 21971 24259
rect 21913 24219 21971 24225
rect 16301 24191 16359 24197
rect 16301 24188 16313 24191
rect 15160 24160 16313 24188
rect 15160 24148 15166 24160
rect 16301 24157 16313 24160
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 17304 24191 17362 24197
rect 17083 24160 17172 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 934 24080 940 24132
rect 992 24120 998 24132
rect 1489 24123 1547 24129
rect 1489 24120 1501 24123
rect 992 24092 1501 24120
rect 992 24080 998 24092
rect 1489 24089 1501 24092
rect 1535 24089 1547 24123
rect 1489 24083 1547 24089
rect 1854 24080 1860 24132
rect 1912 24080 1918 24132
rect 13814 24080 13820 24132
rect 13872 24120 13878 24132
rect 15390 24123 15448 24129
rect 15390 24120 15402 24123
rect 13872 24092 15402 24120
rect 13872 24080 13878 24092
rect 15390 24089 15402 24092
rect 15436 24089 15448 24123
rect 15390 24083 15448 24089
rect 8386 24012 8392 24064
rect 8444 24012 8450 24064
rect 9674 24012 9680 24064
rect 9732 24012 9738 24064
rect 11517 24055 11575 24061
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 12250 24052 12256 24064
rect 11563 24024 12256 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 12250 24012 12256 24024
rect 12308 24012 12314 24064
rect 13722 24012 13728 24064
rect 13780 24052 13786 24064
rect 15286 24052 15292 24064
rect 13780 24024 15292 24052
rect 13780 24012 13786 24024
rect 15286 24012 15292 24024
rect 15344 24012 15350 24064
rect 15746 24012 15752 24064
rect 15804 24012 15810 24064
rect 17144 24052 17172 24160
rect 17304 24157 17316 24191
rect 17350 24157 17362 24191
rect 17304 24151 17362 24157
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 17218 24080 17224 24132
rect 17276 24120 17282 24132
rect 17328 24120 17356 24151
rect 17494 24120 17500 24132
rect 17276 24092 17356 24120
rect 17420 24092 17500 24120
rect 17276 24080 17282 24092
rect 17420 24052 17448 24092
rect 17494 24080 17500 24092
rect 17552 24120 17558 24132
rect 19904 24120 19932 24151
rect 20438 24148 20444 24200
rect 20496 24148 20502 24200
rect 20622 24148 20628 24200
rect 20680 24188 20686 24200
rect 21729 24191 21787 24197
rect 21729 24188 21741 24191
rect 20680 24160 21741 24188
rect 20680 24148 20686 24160
rect 21729 24157 21741 24160
rect 21775 24188 21787 24191
rect 22572 24188 22600 24364
rect 23584 24324 23612 24364
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24394 24392 24400 24404
rect 24075 24364 24400 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 24578 24352 24584 24404
rect 24636 24352 24642 24404
rect 24854 24352 24860 24404
rect 24912 24352 24918 24404
rect 23584 24296 24532 24324
rect 21775 24160 22600 24188
rect 22649 24191 22707 24197
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 22649 24157 22661 24191
rect 22695 24188 22707 24191
rect 23750 24188 23756 24200
rect 22695 24160 23756 24188
rect 22695 24157 22707 24160
rect 22649 24151 22707 24157
rect 19978 24120 19984 24132
rect 17552 24092 19984 24120
rect 17552 24080 17558 24092
rect 19978 24080 19984 24092
rect 20036 24080 20042 24132
rect 20145 24123 20203 24129
rect 20145 24120 20157 24123
rect 20088 24092 20157 24120
rect 17144 24024 17448 24052
rect 19797 24055 19855 24061
rect 19797 24021 19809 24055
rect 19843 24052 19855 24055
rect 20088 24052 20116 24092
rect 20145 24089 20157 24092
rect 20191 24089 20203 24123
rect 20456 24120 20484 24148
rect 22664 24120 22692 24151
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 20456 24092 22692 24120
rect 22916 24123 22974 24129
rect 20145 24083 20203 24089
rect 22916 24089 22928 24123
rect 22962 24089 22974 24123
rect 24504 24120 24532 24296
rect 24596 24188 24624 24352
rect 24872 24324 24900 24352
rect 24872 24296 25360 24324
rect 24670 24216 24676 24268
rect 24728 24256 24734 24268
rect 25332 24265 25360 24296
rect 24949 24259 25007 24265
rect 24949 24256 24961 24259
rect 24728 24228 24961 24256
rect 24728 24216 24734 24228
rect 24949 24225 24961 24228
rect 24995 24225 25007 24259
rect 24949 24219 25007 24225
rect 25317 24259 25375 24265
rect 25317 24225 25329 24259
rect 25363 24225 25375 24259
rect 25317 24219 25375 24225
rect 24765 24191 24823 24197
rect 24765 24188 24777 24191
rect 24596 24160 24777 24188
rect 24765 24157 24777 24160
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 24857 24123 24915 24129
rect 24857 24120 24869 24123
rect 24504 24092 24869 24120
rect 22916 24083 22974 24089
rect 24857 24089 24869 24092
rect 24903 24120 24915 24123
rect 25501 24123 25559 24129
rect 25501 24120 25513 24123
rect 24903 24092 25513 24120
rect 24903 24089 24915 24092
rect 24857 24083 24915 24089
rect 25501 24089 25513 24092
rect 25547 24120 25559 24123
rect 25547 24092 26924 24120
rect 25547 24089 25559 24092
rect 25501 24083 25559 24089
rect 19843 24024 20116 24052
rect 19843 24021 19855 24024
rect 19797 24015 19855 24021
rect 21818 24012 21824 24064
rect 21876 24012 21882 24064
rect 22830 24012 22836 24064
rect 22888 24052 22894 24064
rect 22940 24052 22968 24083
rect 26896 24064 26924 24092
rect 22888 24024 22968 24052
rect 22888 24012 22894 24024
rect 24118 24012 24124 24064
rect 24176 24052 24182 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 24176 24024 24409 24052
rect 24176 24012 24182 24024
rect 24397 24021 24409 24024
rect 24443 24021 24455 24055
rect 24397 24015 24455 24021
rect 25590 24012 25596 24064
rect 25648 24012 25654 24064
rect 25958 24012 25964 24064
rect 26016 24012 26022 24064
rect 26878 24012 26884 24064
rect 26936 24012 26942 24064
rect 1104 23962 31280 23984
rect 1104 23910 4922 23962
rect 4974 23910 4986 23962
rect 5038 23910 5050 23962
rect 5102 23910 5114 23962
rect 5166 23910 5178 23962
rect 5230 23910 5242 23962
rect 5294 23910 10922 23962
rect 10974 23910 10986 23962
rect 11038 23910 11050 23962
rect 11102 23910 11114 23962
rect 11166 23910 11178 23962
rect 11230 23910 11242 23962
rect 11294 23910 16922 23962
rect 16974 23910 16986 23962
rect 17038 23910 17050 23962
rect 17102 23910 17114 23962
rect 17166 23910 17178 23962
rect 17230 23910 17242 23962
rect 17294 23910 22922 23962
rect 22974 23910 22986 23962
rect 23038 23910 23050 23962
rect 23102 23910 23114 23962
rect 23166 23910 23178 23962
rect 23230 23910 23242 23962
rect 23294 23910 28922 23962
rect 28974 23910 28986 23962
rect 29038 23910 29050 23962
rect 29102 23910 29114 23962
rect 29166 23910 29178 23962
rect 29230 23910 29242 23962
rect 29294 23910 31280 23962
rect 1104 23888 31280 23910
rect 8386 23808 8392 23860
rect 8444 23808 8450 23860
rect 8570 23808 8576 23860
rect 8628 23848 8634 23860
rect 9493 23851 9551 23857
rect 9493 23848 9505 23851
rect 8628 23820 9505 23848
rect 8628 23808 8634 23820
rect 9493 23817 9505 23820
rect 9539 23817 9551 23851
rect 9493 23811 9551 23817
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 9861 23851 9919 23857
rect 9861 23848 9873 23851
rect 9732 23820 9873 23848
rect 9732 23808 9738 23820
rect 9861 23817 9873 23820
rect 9907 23817 9919 23851
rect 9861 23811 9919 23817
rect 13446 23808 13452 23860
rect 13504 23848 13510 23860
rect 13722 23848 13728 23860
rect 13504 23820 13728 23848
rect 13504 23808 13510 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 13814 23808 13820 23860
rect 13872 23808 13878 23860
rect 13909 23851 13967 23857
rect 13909 23817 13921 23851
rect 13955 23817 13967 23851
rect 13909 23811 13967 23817
rect 14277 23851 14335 23857
rect 14277 23817 14289 23851
rect 14323 23848 14335 23851
rect 14366 23848 14372 23860
rect 14323 23820 14372 23848
rect 14323 23817 14335 23820
rect 14277 23811 14335 23817
rect 8288 23783 8346 23789
rect 8288 23749 8300 23783
rect 8334 23780 8346 23783
rect 8404 23780 8432 23808
rect 8334 23752 8432 23780
rect 12820 23752 13584 23780
rect 8334 23749 8346 23752
rect 8288 23743 8346 23749
rect 12820 23724 12848 23752
rect 13556 23724 13584 23752
rect 4985 23715 5043 23721
rect 4985 23681 4997 23715
rect 5031 23712 5043 23715
rect 5445 23715 5503 23721
rect 5445 23712 5457 23715
rect 5031 23684 5457 23712
rect 5031 23681 5043 23684
rect 4985 23675 5043 23681
rect 5445 23681 5457 23684
rect 5491 23681 5503 23715
rect 5445 23675 5503 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23712 8079 23715
rect 8110 23712 8116 23724
rect 8067 23684 8116 23712
rect 8067 23681 8079 23684
rect 8021 23675 8079 23681
rect 8110 23672 8116 23684
rect 8168 23672 8174 23724
rect 9950 23672 9956 23724
rect 10008 23712 10014 23724
rect 10008 23684 12434 23712
rect 10008 23672 10014 23684
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23613 5135 23647
rect 5077 23607 5135 23613
rect 5261 23647 5319 23653
rect 5261 23613 5273 23647
rect 5307 23644 5319 23647
rect 5350 23644 5356 23656
rect 5307 23616 5356 23644
rect 5307 23613 5319 23616
rect 5261 23607 5319 23613
rect 4614 23468 4620 23520
rect 4672 23468 4678 23520
rect 5092 23508 5120 23607
rect 5350 23604 5356 23616
rect 5408 23644 5414 23656
rect 5902 23644 5908 23656
rect 5408 23616 5908 23644
rect 5408 23604 5414 23616
rect 5902 23604 5908 23616
rect 5960 23604 5966 23656
rect 5994 23604 6000 23656
rect 6052 23604 6058 23656
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10045 23647 10103 23653
rect 10045 23644 10057 23647
rect 9916 23616 10057 23644
rect 9916 23604 9922 23616
rect 10045 23613 10057 23616
rect 10091 23613 10103 23647
rect 10045 23607 10103 23613
rect 9401 23579 9459 23585
rect 9401 23545 9413 23579
rect 9447 23576 9459 23579
rect 10778 23576 10784 23588
rect 9447 23548 10784 23576
rect 9447 23545 9459 23548
rect 9401 23539 9459 23545
rect 10778 23536 10784 23548
rect 10836 23536 10842 23588
rect 12406 23576 12434 23684
rect 12802 23672 12808 23724
rect 12860 23672 12866 23724
rect 12989 23715 13047 23721
rect 12989 23681 13001 23715
rect 13035 23681 13047 23715
rect 12989 23675 13047 23681
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13446 23712 13452 23724
rect 13127 23684 13452 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 13004 23644 13032 23675
rect 13446 23672 13452 23684
rect 13504 23672 13510 23724
rect 13538 23672 13544 23724
rect 13596 23672 13602 23724
rect 13633 23715 13691 23721
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13924 23712 13952 23811
rect 14366 23808 14372 23820
rect 14424 23808 14430 23860
rect 14737 23851 14795 23857
rect 14737 23817 14749 23851
rect 14783 23848 14795 23851
rect 15102 23848 15108 23860
rect 14783 23820 15108 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 15102 23808 15108 23820
rect 15160 23808 15166 23860
rect 16114 23808 16120 23860
rect 16172 23808 16178 23860
rect 17586 23808 17592 23860
rect 17644 23808 17650 23860
rect 18322 23808 18328 23860
rect 18380 23808 18386 23860
rect 20254 23808 20260 23860
rect 20312 23808 20318 23860
rect 21174 23808 21180 23860
rect 21232 23808 21238 23860
rect 21818 23808 21824 23860
rect 21876 23808 21882 23860
rect 23477 23851 23535 23857
rect 23477 23817 23489 23851
rect 23523 23848 23535 23851
rect 23842 23848 23848 23860
rect 23523 23820 23848 23848
rect 23523 23817 23535 23820
rect 23477 23811 23535 23817
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24118 23808 24124 23860
rect 24176 23808 24182 23860
rect 24213 23851 24271 23857
rect 24213 23817 24225 23851
rect 24259 23817 24271 23851
rect 24213 23811 24271 23817
rect 16132 23721 16160 23808
rect 17862 23780 17868 23792
rect 17236 23752 17868 23780
rect 17236 23724 17264 23752
rect 17862 23740 17868 23752
rect 17920 23740 17926 23792
rect 13679 23684 13952 23712
rect 15861 23715 15919 23721
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 15861 23681 15873 23715
rect 15907 23712 15919 23715
rect 16117 23715 16175 23721
rect 15907 23684 16068 23712
rect 15907 23681 15919 23684
rect 15861 23675 15919 23681
rect 13906 23644 13912 23656
rect 13004 23616 13912 23644
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 14369 23647 14427 23653
rect 14369 23613 14381 23647
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 13446 23576 13452 23588
rect 12406 23548 13452 23576
rect 13446 23536 13452 23548
rect 13504 23576 13510 23588
rect 14384 23576 14412 23607
rect 14550 23604 14556 23656
rect 14608 23604 14614 23656
rect 16040 23644 16068 23684
rect 16117 23681 16129 23715
rect 16163 23681 16175 23715
rect 16117 23675 16175 23681
rect 16206 23672 16212 23724
rect 16264 23712 16270 23724
rect 16393 23715 16451 23721
rect 16393 23712 16405 23715
rect 16264 23684 16405 23712
rect 16264 23672 16270 23684
rect 16393 23681 16405 23684
rect 16439 23681 16451 23715
rect 16393 23675 16451 23681
rect 17218 23672 17224 23724
rect 17276 23672 17282 23724
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23712 17463 23715
rect 18340 23712 18368 23808
rect 17451 23684 18368 23712
rect 18693 23715 18751 23721
rect 17451 23681 17463 23684
rect 17405 23675 17463 23681
rect 18693 23681 18705 23715
rect 18739 23712 18751 23715
rect 19978 23712 19984 23724
rect 18739 23684 19984 23712
rect 18739 23681 18751 23684
rect 18693 23675 18751 23681
rect 19978 23672 19984 23684
rect 20036 23712 20042 23724
rect 20073 23715 20131 23721
rect 20073 23712 20085 23715
rect 20036 23684 20085 23712
rect 20036 23672 20042 23684
rect 20073 23681 20085 23684
rect 20119 23681 20131 23715
rect 20272 23712 20300 23808
rect 20340 23783 20398 23789
rect 20340 23749 20352 23783
rect 20386 23780 20398 23783
rect 21192 23780 21220 23808
rect 20386 23752 21220 23780
rect 22557 23783 22615 23789
rect 20386 23749 20398 23752
rect 20340 23743 20398 23749
rect 22557 23749 22569 23783
rect 22603 23780 22615 23783
rect 22646 23780 22652 23792
rect 22603 23752 22652 23780
rect 22603 23749 22615 23752
rect 22557 23743 22615 23749
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 23750 23740 23756 23792
rect 23808 23780 23814 23792
rect 23808 23752 23980 23780
rect 23808 23740 23814 23752
rect 22833 23715 22891 23721
rect 20272 23684 21220 23712
rect 20073 23675 20131 23681
rect 16040 23616 16252 23644
rect 13504 23548 14412 23576
rect 13504 23536 13510 23548
rect 9214 23508 9220 23520
rect 5092 23480 9220 23508
rect 9214 23468 9220 23480
rect 9272 23468 9278 23520
rect 9766 23468 9772 23520
rect 9824 23508 9830 23520
rect 10594 23508 10600 23520
rect 9824 23480 10600 23508
rect 9824 23468 9830 23480
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12621 23511 12679 23517
rect 12621 23508 12633 23511
rect 12492 23480 12633 23508
rect 12492 23468 12498 23480
rect 12621 23477 12633 23480
rect 12667 23477 12679 23511
rect 14568 23508 14596 23604
rect 16224 23585 16252 23616
rect 16209 23579 16267 23585
rect 16209 23545 16221 23579
rect 16255 23545 16267 23579
rect 16209 23539 16267 23545
rect 18874 23508 18880 23520
rect 14568 23480 18880 23508
rect 12621 23471 12679 23477
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 20254 23468 20260 23520
rect 20312 23508 20318 23520
rect 20990 23508 20996 23520
rect 20312 23480 20996 23508
rect 20312 23468 20318 23480
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21192 23508 21220 23684
rect 22833 23681 22845 23715
rect 22879 23712 22891 23715
rect 23474 23712 23480 23724
rect 22879 23684 23480 23712
rect 22879 23681 22891 23684
rect 22833 23675 22891 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 23566 23672 23572 23724
rect 23624 23712 23630 23724
rect 23624 23684 23888 23712
rect 23624 23672 23630 23684
rect 23860 23656 23888 23684
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 22066 23616 22385 23644
rect 22066 23588 22094 23616
rect 22373 23613 22385 23616
rect 22419 23613 22431 23647
rect 22373 23607 22431 23613
rect 22741 23647 22799 23653
rect 22741 23613 22753 23647
rect 22787 23613 22799 23647
rect 22741 23607 22799 23613
rect 21453 23579 21511 23585
rect 21453 23545 21465 23579
rect 21499 23576 21511 23579
rect 22066 23576 22100 23588
rect 21499 23548 22100 23576
rect 21499 23545 21511 23548
rect 21453 23539 21511 23545
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 22756 23576 22784 23607
rect 23658 23604 23664 23656
rect 23716 23604 23722 23656
rect 23842 23604 23848 23656
rect 23900 23604 23906 23656
rect 23952 23644 23980 23752
rect 24029 23715 24087 23721
rect 24029 23681 24041 23715
rect 24075 23712 24087 23715
rect 24136 23712 24164 23808
rect 24228 23780 24256 23811
rect 25590 23808 25596 23860
rect 25648 23848 25654 23860
rect 25777 23851 25835 23857
rect 25777 23848 25789 23851
rect 25648 23820 25789 23848
rect 25648 23808 25654 23820
rect 25777 23817 25789 23820
rect 25823 23817 25835 23851
rect 25777 23811 25835 23817
rect 25958 23808 25964 23860
rect 26016 23808 26022 23860
rect 24550 23783 24608 23789
rect 24550 23780 24562 23783
rect 24228 23752 24562 23780
rect 24550 23749 24562 23752
rect 24596 23749 24608 23783
rect 24550 23743 24608 23749
rect 24075 23684 24164 23712
rect 25976 23712 26004 23808
rect 26697 23715 26755 23721
rect 26697 23712 26709 23715
rect 25976 23684 26709 23712
rect 24075 23681 24087 23684
rect 24029 23675 24087 23681
rect 26697 23681 26709 23684
rect 26743 23681 26755 23715
rect 26697 23675 26755 23681
rect 24118 23644 24124 23656
rect 23952 23616 24124 23644
rect 24118 23604 24124 23616
rect 24176 23644 24182 23656
rect 24305 23647 24363 23653
rect 24305 23644 24317 23647
rect 24176 23616 24317 23644
rect 24176 23604 24182 23616
rect 24305 23613 24317 23616
rect 24351 23613 24363 23647
rect 24305 23607 24363 23613
rect 26326 23604 26332 23656
rect 26384 23604 26390 23656
rect 22756 23548 23336 23576
rect 22557 23511 22615 23517
rect 22557 23508 22569 23511
rect 21192 23480 22569 23508
rect 22557 23477 22569 23480
rect 22603 23477 22615 23511
rect 22557 23471 22615 23477
rect 23014 23468 23020 23520
rect 23072 23468 23078 23520
rect 23106 23468 23112 23520
rect 23164 23468 23170 23520
rect 23308 23508 23336 23548
rect 23750 23508 23756 23520
rect 23308 23480 23756 23508
rect 23750 23468 23756 23480
rect 23808 23468 23814 23520
rect 25222 23468 25228 23520
rect 25280 23508 25286 23520
rect 25685 23511 25743 23517
rect 25685 23508 25697 23511
rect 25280 23480 25697 23508
rect 25280 23468 25286 23480
rect 25685 23477 25697 23480
rect 25731 23477 25743 23511
rect 25685 23471 25743 23477
rect 26510 23468 26516 23520
rect 26568 23468 26574 23520
rect 1104 23418 31280 23440
rect 1104 23366 4182 23418
rect 4234 23366 4246 23418
rect 4298 23366 4310 23418
rect 4362 23366 4374 23418
rect 4426 23366 4438 23418
rect 4490 23366 4502 23418
rect 4554 23366 10182 23418
rect 10234 23366 10246 23418
rect 10298 23366 10310 23418
rect 10362 23366 10374 23418
rect 10426 23366 10438 23418
rect 10490 23366 10502 23418
rect 10554 23366 16182 23418
rect 16234 23366 16246 23418
rect 16298 23366 16310 23418
rect 16362 23366 16374 23418
rect 16426 23366 16438 23418
rect 16490 23366 16502 23418
rect 16554 23366 22182 23418
rect 22234 23366 22246 23418
rect 22298 23366 22310 23418
rect 22362 23366 22374 23418
rect 22426 23366 22438 23418
rect 22490 23366 22502 23418
rect 22554 23366 28182 23418
rect 28234 23366 28246 23418
rect 28298 23366 28310 23418
rect 28362 23366 28374 23418
rect 28426 23366 28438 23418
rect 28490 23366 28502 23418
rect 28554 23366 31280 23418
rect 1104 23344 31280 23366
rect 4706 23264 4712 23316
rect 4764 23264 4770 23316
rect 7006 23304 7012 23316
rect 6656 23276 7012 23304
rect 4724 23168 4752 23264
rect 4801 23171 4859 23177
rect 4801 23168 4813 23171
rect 4724 23140 4813 23168
rect 4801 23137 4813 23140
rect 4847 23137 4859 23171
rect 4801 23131 4859 23137
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23100 4491 23103
rect 4614 23100 4620 23112
rect 4479 23072 4620 23100
rect 4479 23069 4491 23072
rect 4433 23063 4491 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6656 23109 6684 23276
rect 7006 23264 7012 23276
rect 7064 23304 7070 23316
rect 9950 23304 9956 23316
rect 7064 23276 9956 23304
rect 7064 23264 7070 23276
rect 9950 23264 9956 23276
rect 10008 23264 10014 23316
rect 10870 23264 10876 23316
rect 10928 23304 10934 23316
rect 11514 23304 11520 23316
rect 10928 23276 11520 23304
rect 10928 23264 10934 23276
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 11793 23307 11851 23313
rect 11793 23273 11805 23307
rect 11839 23273 11851 23307
rect 11793 23267 11851 23273
rect 8757 23239 8815 23245
rect 8757 23205 8769 23239
rect 8803 23236 8815 23239
rect 11808 23236 11836 23267
rect 13906 23264 13912 23316
rect 13964 23264 13970 23316
rect 15749 23307 15807 23313
rect 15749 23273 15761 23307
rect 15795 23304 15807 23307
rect 16022 23304 16028 23316
rect 15795 23276 16028 23304
rect 15795 23273 15807 23276
rect 15749 23267 15807 23273
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 22373 23307 22431 23313
rect 22373 23273 22385 23307
rect 22419 23304 22431 23307
rect 22646 23304 22652 23316
rect 22419 23276 22652 23304
rect 22419 23273 22431 23276
rect 22373 23267 22431 23273
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22888 23276 22937 23304
rect 22888 23264 22894 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 22925 23267 22983 23273
rect 23474 23264 23480 23316
rect 23532 23304 23538 23316
rect 23661 23307 23719 23313
rect 23661 23304 23673 23307
rect 23532 23276 23673 23304
rect 23532 23264 23538 23276
rect 23661 23273 23673 23276
rect 23707 23273 23719 23307
rect 23661 23267 23719 23273
rect 24486 23264 24492 23316
rect 24544 23304 24550 23316
rect 26326 23304 26332 23316
rect 24544 23276 26332 23304
rect 24544 23264 24550 23276
rect 26326 23264 26332 23276
rect 26384 23264 26390 23316
rect 11882 23236 11888 23248
rect 8803 23208 10364 23236
rect 11808 23208 11888 23236
rect 8803 23205 8815 23208
rect 8757 23199 8815 23205
rect 6822 23128 6828 23180
rect 6880 23128 6886 23180
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9401 23171 9459 23177
rect 9401 23168 9413 23171
rect 9272 23140 9413 23168
rect 9272 23128 9278 23140
rect 9401 23137 9413 23140
rect 9447 23137 9459 23171
rect 9401 23131 9459 23137
rect 9585 23171 9643 23177
rect 9585 23137 9597 23171
rect 9631 23168 9643 23171
rect 9766 23168 9772 23180
rect 9631 23140 9772 23168
rect 9631 23137 9643 23140
rect 9585 23131 9643 23137
rect 6641 23103 6699 23109
rect 6641 23069 6653 23103
rect 6687 23069 6699 23103
rect 6641 23063 6699 23069
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 8110 23100 8116 23112
rect 7423 23072 8116 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 8110 23060 8116 23072
rect 8168 23060 8174 23112
rect 9416 23100 9444 23131
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 10336 23177 10364 23208
rect 11882 23196 11888 23208
rect 11940 23196 11946 23248
rect 10321 23171 10379 23177
rect 10321 23137 10333 23171
rect 10367 23168 10379 23171
rect 11698 23168 11704 23180
rect 10367 23140 10548 23168
rect 10367 23137 10379 23140
rect 10321 23131 10379 23137
rect 9858 23100 9864 23112
rect 9416 23072 9864 23100
rect 9858 23060 9864 23072
rect 9916 23100 9922 23112
rect 10226 23100 10232 23112
rect 9916 23072 10232 23100
rect 9916 23060 9922 23072
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 10520 23109 10548 23140
rect 10704 23140 11704 23168
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 10704 23109 10732 23140
rect 11698 23128 11704 23140
rect 11756 23128 11762 23180
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23168 11851 23171
rect 12434 23168 12440 23180
rect 11839 23140 12440 23168
rect 11839 23137 11851 23140
rect 11793 23131 11851 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 12526 23128 12532 23180
rect 12584 23128 12590 23180
rect 13924 23168 13952 23264
rect 14645 23171 14703 23177
rect 14645 23168 14657 23171
rect 13924 23140 14657 23168
rect 14645 23137 14657 23140
rect 14691 23137 14703 23171
rect 14645 23131 14703 23137
rect 15197 23171 15255 23177
rect 15197 23137 15209 23171
rect 15243 23168 15255 23171
rect 15470 23168 15476 23180
rect 15243 23140 15476 23168
rect 15243 23137 15255 23140
rect 15197 23131 15255 23137
rect 15470 23128 15476 23140
rect 15528 23168 15534 23180
rect 17770 23168 17776 23180
rect 15528 23140 17776 23168
rect 15528 23128 15534 23140
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 20438 23128 20444 23180
rect 20496 23168 20502 23180
rect 21177 23171 21235 23177
rect 21177 23168 21189 23171
rect 20496 23140 21189 23168
rect 20496 23128 20502 23140
rect 21177 23137 21189 23140
rect 21223 23137 21235 23171
rect 21177 23131 21235 23137
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 24176 23140 24532 23168
rect 24176 23128 24182 23140
rect 10689 23103 10747 23109
rect 10689 23100 10701 23103
rect 10652 23072 10701 23100
rect 10652 23060 10658 23072
rect 10689 23069 10701 23072
rect 10735 23069 10747 23103
rect 10689 23063 10747 23069
rect 10778 23060 10784 23112
rect 10836 23060 10842 23112
rect 10870 23060 10876 23112
rect 10928 23060 10934 23112
rect 11885 23103 11943 23109
rect 11885 23076 11897 23103
rect 11808 23069 11897 23076
rect 11931 23069 11943 23103
rect 11808 23063 11943 23069
rect 11808 23048 11921 23063
rect 12250 23060 12256 23112
rect 12308 23060 12314 23112
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 15289 23103 15347 23109
rect 15289 23100 15301 23103
rect 12676 23072 15301 23100
rect 12676 23060 12682 23072
rect 15289 23069 15301 23072
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 15746 23100 15752 23112
rect 15427 23072 15752 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 19334 23060 19340 23112
rect 19392 23060 19398 23112
rect 21266 23060 21272 23112
rect 21324 23100 21330 23112
rect 21821 23103 21879 23109
rect 21821 23100 21833 23103
rect 21324 23072 21833 23100
rect 21324 23060 21330 23072
rect 21821 23069 21833 23072
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22094 23060 22100 23112
rect 22152 23060 22158 23112
rect 22189 23103 22247 23109
rect 22189 23069 22201 23103
rect 22235 23100 22247 23103
rect 22646 23100 22652 23112
rect 22235 23072 22652 23100
rect 22235 23069 22247 23072
rect 22189 23063 22247 23069
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 23937 23103 23995 23109
rect 23937 23069 23949 23103
rect 23983 23100 23995 23103
rect 24213 23103 24271 23109
rect 23983 23072 24164 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 5068 23035 5126 23041
rect 5068 23001 5080 23035
rect 5114 23032 5126 23035
rect 5350 23032 5356 23044
rect 5114 23004 5356 23032
rect 5114 23001 5126 23004
rect 5068 22995 5126 23001
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 7644 23035 7702 23041
rect 7644 23001 7656 23035
rect 7690 23032 7702 23035
rect 7742 23032 7748 23044
rect 7690 23004 7748 23032
rect 7690 23001 7702 23004
rect 7644 22995 7702 23001
rect 7742 22992 7748 23004
rect 7800 22992 7806 23044
rect 9309 23035 9367 23041
rect 9309 23001 9321 23035
rect 9355 23032 9367 23035
rect 9769 23035 9827 23041
rect 9769 23032 9781 23035
rect 9355 23004 9781 23032
rect 9355 23001 9367 23004
rect 9309 22995 9367 23001
rect 9769 23001 9781 23004
rect 9815 23001 9827 23035
rect 9769 22995 9827 23001
rect 11606 22992 11612 23044
rect 11664 22992 11670 23044
rect 4246 22924 4252 22976
rect 4304 22924 4310 22976
rect 6178 22924 6184 22976
rect 6236 22924 6242 22976
rect 6270 22924 6276 22976
rect 6328 22924 6334 22976
rect 6730 22924 6736 22976
rect 6788 22924 6794 22976
rect 8938 22924 8944 22976
rect 8996 22924 9002 22976
rect 11057 22967 11115 22973
rect 11057 22933 11069 22967
rect 11103 22964 11115 22967
rect 11808 22964 11836 23048
rect 12774 23035 12832 23041
rect 12774 23032 12786 23035
rect 12452 23004 12786 23032
rect 11103 22936 11836 22964
rect 11103 22933 11115 22936
rect 11057 22927 11115 22933
rect 12066 22924 12072 22976
rect 12124 22924 12130 22976
rect 12452 22973 12480 23004
rect 12774 23001 12786 23004
rect 12820 23001 12832 23035
rect 19352 23032 19380 23060
rect 20441 23035 20499 23041
rect 20441 23032 20453 23035
rect 19352 23004 20453 23032
rect 12774 22995 12832 23001
rect 20441 23001 20453 23004
rect 20487 23001 20499 23035
rect 22005 23035 22063 23041
rect 22005 23032 22017 23035
rect 20441 22995 20499 23001
rect 21836 23004 22017 23032
rect 21836 22976 21864 23004
rect 22005 23001 22017 23004
rect 22051 23001 22063 23035
rect 22664 23032 22692 23060
rect 23290 23032 23296 23044
rect 22664 23004 23296 23032
rect 22005 22995 22063 23001
rect 23290 22992 23296 23004
rect 23348 22992 23354 23044
rect 12437 22967 12495 22973
rect 12437 22933 12449 22967
rect 12483 22933 12495 22967
rect 12437 22927 12495 22933
rect 14090 22924 14096 22976
rect 14148 22924 14154 22976
rect 21818 22924 21824 22976
rect 21876 22924 21882 22976
rect 23860 22964 23888 23063
rect 24026 22992 24032 23044
rect 24084 22992 24090 23044
rect 24136 23032 24164 23072
rect 24213 23069 24225 23103
rect 24259 23100 24271 23103
rect 24394 23100 24400 23112
rect 24259 23072 24400 23100
rect 24259 23069 24271 23072
rect 24213 23063 24271 23069
rect 24394 23060 24400 23072
rect 24452 23060 24458 23112
rect 24504 23100 24532 23140
rect 25038 23100 25044 23112
rect 24504 23072 25044 23100
rect 25038 23060 25044 23072
rect 25096 23100 25102 23112
rect 25869 23103 25927 23109
rect 25869 23100 25881 23103
rect 25096 23072 25881 23100
rect 25096 23060 25102 23072
rect 25869 23069 25881 23072
rect 25915 23069 25927 23103
rect 25869 23063 25927 23069
rect 26510 23060 26516 23112
rect 26568 23060 26574 23112
rect 25222 23032 25228 23044
rect 24136 23004 25228 23032
rect 25222 22992 25228 23004
rect 25280 22992 25286 23044
rect 25624 23035 25682 23041
rect 25624 23001 25636 23035
rect 25670 23032 25682 23035
rect 26528 23032 26556 23060
rect 25670 23004 26556 23032
rect 25670 23001 25682 23004
rect 25624 22995 25682 23001
rect 24394 22964 24400 22976
rect 23860 22936 24400 22964
rect 24394 22924 24400 22936
rect 24452 22924 24458 22976
rect 1104 22874 31280 22896
rect 1104 22822 4922 22874
rect 4974 22822 4986 22874
rect 5038 22822 5050 22874
rect 5102 22822 5114 22874
rect 5166 22822 5178 22874
rect 5230 22822 5242 22874
rect 5294 22822 10922 22874
rect 10974 22822 10986 22874
rect 11038 22822 11050 22874
rect 11102 22822 11114 22874
rect 11166 22822 11178 22874
rect 11230 22822 11242 22874
rect 11294 22822 16922 22874
rect 16974 22822 16986 22874
rect 17038 22822 17050 22874
rect 17102 22822 17114 22874
rect 17166 22822 17178 22874
rect 17230 22822 17242 22874
rect 17294 22822 22922 22874
rect 22974 22822 22986 22874
rect 23038 22822 23050 22874
rect 23102 22822 23114 22874
rect 23166 22822 23178 22874
rect 23230 22822 23242 22874
rect 23294 22822 28922 22874
rect 28974 22822 28986 22874
rect 29038 22822 29050 22874
rect 29102 22822 29114 22874
rect 29166 22822 29178 22874
rect 29230 22822 29242 22874
rect 29294 22822 31280 22874
rect 1104 22800 31280 22822
rect 4246 22720 4252 22772
rect 4304 22720 4310 22772
rect 5350 22720 5356 22772
rect 5408 22720 5414 22772
rect 6270 22720 6276 22772
rect 6328 22720 6334 22772
rect 6457 22763 6515 22769
rect 6457 22729 6469 22763
rect 6503 22760 6515 22763
rect 6730 22760 6736 22772
rect 6503 22732 6736 22760
rect 6503 22729 6515 22732
rect 6457 22723 6515 22729
rect 6730 22720 6736 22732
rect 6788 22720 6794 22772
rect 7190 22720 7196 22772
rect 7248 22720 7254 22772
rect 7742 22720 7748 22772
rect 7800 22760 7806 22772
rect 7837 22763 7895 22769
rect 7837 22760 7849 22763
rect 7800 22732 7849 22760
rect 7800 22720 7806 22732
rect 7837 22729 7849 22732
rect 7883 22729 7895 22763
rect 7837 22723 7895 22729
rect 8938 22720 8944 22772
rect 8996 22720 9002 22772
rect 11606 22720 11612 22772
rect 11664 22720 11670 22772
rect 12250 22720 12256 22772
rect 12308 22760 12314 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12308 22732 13001 22760
rect 12308 22720 12314 22732
rect 12989 22729 13001 22732
rect 13035 22729 13047 22763
rect 12989 22723 13047 22729
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 14090 22760 14096 22772
rect 13403 22732 14096 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 14369 22763 14427 22769
rect 14369 22729 14381 22763
rect 14415 22729 14427 22763
rect 14918 22760 14924 22772
rect 14369 22723 14427 22729
rect 14660 22732 14924 22760
rect 4148 22695 4206 22701
rect 4148 22661 4160 22695
rect 4194 22692 4206 22695
rect 4264 22692 4292 22720
rect 4194 22664 4292 22692
rect 4194 22661 4206 22664
rect 4148 22655 4206 22661
rect 5537 22627 5595 22633
rect 5537 22593 5549 22627
rect 5583 22624 5595 22627
rect 6288 22624 6316 22720
rect 7208 22692 7236 22720
rect 7377 22695 7435 22701
rect 7377 22692 7389 22695
rect 7208 22664 7389 22692
rect 7377 22661 7389 22664
rect 7423 22661 7435 22695
rect 7377 22655 7435 22661
rect 5583 22596 6316 22624
rect 5583 22593 5595 22596
rect 5537 22587 5595 22593
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 7193 22627 7251 22633
rect 7193 22624 7205 22627
rect 6420 22596 7205 22624
rect 6420 22584 6426 22596
rect 7193 22593 7205 22596
rect 7239 22593 7251 22627
rect 7193 22587 7251 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22593 7527 22627
rect 7469 22587 7527 22593
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22624 7619 22627
rect 7650 22624 7656 22636
rect 7607 22596 7656 22624
rect 7607 22593 7619 22596
rect 7561 22587 7619 22593
rect 3878 22516 3884 22568
rect 3936 22516 3942 22568
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 7009 22559 7067 22565
rect 7009 22556 7021 22559
rect 6236 22528 7021 22556
rect 6236 22516 6242 22528
rect 7009 22525 7021 22528
rect 7055 22556 7067 22559
rect 7484 22556 7512 22587
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 8021 22627 8079 22633
rect 8021 22593 8033 22627
rect 8067 22624 8079 22627
rect 8956 22624 8984 22720
rect 8067 22596 8984 22624
rect 8067 22593 8079 22596
rect 8021 22587 8079 22593
rect 7055 22528 7512 22556
rect 7055 22525 7067 22528
rect 7009 22519 7067 22525
rect 5261 22491 5319 22497
rect 5261 22457 5273 22491
rect 5307 22488 5319 22491
rect 5994 22488 6000 22500
rect 5307 22460 6000 22488
rect 5307 22457 5319 22460
rect 5261 22451 5319 22457
rect 5994 22448 6000 22460
rect 6052 22488 6058 22500
rect 6362 22488 6368 22500
rect 6052 22460 6368 22488
rect 6052 22448 6058 22460
rect 6362 22448 6368 22460
rect 6420 22448 6426 22500
rect 7745 22491 7803 22497
rect 7745 22457 7757 22491
rect 7791 22488 7803 22491
rect 11624 22488 11652 22720
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 14384 22692 14412 22723
rect 14660 22701 14688 22732
rect 14918 22720 14924 22732
rect 14976 22720 14982 22772
rect 23750 22720 23756 22772
rect 23808 22720 23814 22772
rect 24121 22763 24179 22769
rect 24121 22729 24133 22763
rect 24167 22760 24179 22763
rect 24486 22760 24492 22772
rect 24167 22732 24492 22760
rect 24167 22729 24179 22732
rect 24121 22723 24179 22729
rect 24486 22720 24492 22732
rect 24544 22720 24550 22772
rect 11940 22664 14412 22692
rect 14645 22695 14703 22701
rect 11940 22652 11946 22664
rect 14645 22661 14657 22695
rect 14691 22661 14703 22695
rect 14645 22655 14703 22661
rect 14734 22652 14740 22704
rect 14792 22652 14798 22704
rect 23952 22664 24808 22692
rect 23952 22636 23980 22664
rect 24780 22636 24808 22664
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 14458 22584 14464 22636
rect 14516 22624 14522 22636
rect 14553 22627 14611 22633
rect 14553 22624 14565 22627
rect 14516 22596 14565 22624
rect 14516 22584 14522 22596
rect 14553 22593 14565 22596
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 14921 22627 14979 22633
rect 14921 22593 14933 22627
rect 14967 22624 14979 22627
rect 15102 22624 15108 22636
rect 14967 22596 15108 22624
rect 14967 22593 14979 22596
rect 14921 22587 14979 22593
rect 15102 22584 15108 22596
rect 15160 22584 15166 22636
rect 23934 22584 23940 22636
rect 23992 22584 23998 22636
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 13633 22559 13691 22565
rect 13633 22525 13645 22559
rect 13679 22556 13691 22559
rect 13722 22556 13728 22568
rect 13679 22528 13728 22556
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 13722 22516 13728 22528
rect 13780 22556 13786 22568
rect 15194 22556 15200 22568
rect 13780 22528 15200 22556
rect 13780 22516 13786 22528
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 24118 22516 24124 22568
rect 24176 22556 24182 22568
rect 24228 22556 24256 22587
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 24176 22528 24256 22556
rect 24176 22516 24182 22528
rect 7791 22460 11652 22488
rect 7791 22457 7803 22460
rect 7745 22451 7803 22457
rect 12894 22448 12900 22500
rect 12952 22488 12958 22500
rect 16758 22488 16764 22500
rect 12952 22460 16764 22488
rect 12952 22448 12958 22460
rect 16758 22448 16764 22460
rect 16816 22488 16822 22500
rect 23658 22488 23664 22500
rect 16816 22460 23664 22488
rect 16816 22448 16822 22460
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 18322 22420 18328 22432
rect 17000 22392 18328 22420
rect 17000 22380 17006 22392
rect 18322 22380 18328 22392
rect 18380 22380 18386 22432
rect 1104 22330 31280 22352
rect 1104 22278 4182 22330
rect 4234 22278 4246 22330
rect 4298 22278 4310 22330
rect 4362 22278 4374 22330
rect 4426 22278 4438 22330
rect 4490 22278 4502 22330
rect 4554 22278 10182 22330
rect 10234 22278 10246 22330
rect 10298 22278 10310 22330
rect 10362 22278 10374 22330
rect 10426 22278 10438 22330
rect 10490 22278 10502 22330
rect 10554 22278 16182 22330
rect 16234 22278 16246 22330
rect 16298 22278 16310 22330
rect 16362 22278 16374 22330
rect 16426 22278 16438 22330
rect 16490 22278 16502 22330
rect 16554 22278 22182 22330
rect 22234 22278 22246 22330
rect 22298 22278 22310 22330
rect 22362 22278 22374 22330
rect 22426 22278 22438 22330
rect 22490 22278 22502 22330
rect 22554 22278 28182 22330
rect 28234 22278 28246 22330
rect 28298 22278 28310 22330
rect 28362 22278 28374 22330
rect 28426 22278 28438 22330
rect 28490 22278 28502 22330
rect 28554 22278 31280 22330
rect 1104 22256 31280 22278
rect 9766 22216 9772 22228
rect 9646 22188 9772 22216
rect 9646 22148 9674 22188
rect 9766 22176 9772 22188
rect 9824 22216 9830 22228
rect 9824 22188 12940 22216
rect 9824 22176 9830 22188
rect 12912 22160 12940 22188
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 15470 22216 15476 22228
rect 15252 22188 15476 22216
rect 15252 22176 15258 22188
rect 15470 22176 15476 22188
rect 15528 22176 15534 22228
rect 16592 22188 19012 22216
rect 16592 22160 16620 22188
rect 8496 22120 9674 22148
rect 5718 22040 5724 22092
rect 5776 22080 5782 22092
rect 8110 22080 8116 22092
rect 5776 22052 8116 22080
rect 5776 22040 5782 22052
rect 8110 22040 8116 22052
rect 8168 22080 8174 22092
rect 8496 22089 8524 22120
rect 10778 22108 10784 22160
rect 10836 22148 10842 22160
rect 11514 22148 11520 22160
rect 10836 22120 11520 22148
rect 10836 22108 10842 22120
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 12894 22108 12900 22160
rect 12952 22108 12958 22160
rect 14090 22108 14096 22160
rect 14148 22108 14154 22160
rect 16574 22108 16580 22160
rect 16632 22108 16638 22160
rect 17586 22148 17592 22160
rect 17420 22120 17592 22148
rect 8297 22083 8355 22089
rect 8297 22080 8309 22083
rect 8168 22052 8309 22080
rect 8168 22040 8174 22052
rect 8297 22049 8309 22052
rect 8343 22049 8355 22083
rect 8297 22043 8355 22049
rect 8481 22083 8539 22089
rect 8481 22049 8493 22083
rect 8527 22080 8539 22083
rect 13262 22080 13268 22092
rect 8527 22052 8561 22080
rect 8680 22052 13268 22080
rect 8527 22049 8539 22052
rect 8481 22043 8539 22049
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 8680 22012 8708 22052
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 17420 22089 17448 22120
rect 17586 22108 17592 22120
rect 17644 22108 17650 22160
rect 17405 22083 17463 22089
rect 17405 22049 17417 22083
rect 17451 22049 17463 22083
rect 17405 22043 17463 22049
rect 17957 22083 18015 22089
rect 17957 22049 17969 22083
rect 18003 22080 18015 22083
rect 18874 22080 18880 22092
rect 18003 22052 18880 22080
rect 18003 22049 18015 22052
rect 17957 22043 18015 22049
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 7432 21984 8708 22012
rect 7432 21972 7438 21984
rect 9306 21972 9312 22024
rect 9364 21972 9370 22024
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 22012 11115 22015
rect 11103 21984 11652 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 11624 21888 11652 21984
rect 13078 21972 13084 22024
rect 13136 22012 13142 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 13136 21984 14657 22012
rect 13136 21972 13142 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 15565 22015 15623 22021
rect 14645 21975 14703 21981
rect 14752 21984 15516 22012
rect 11974 21904 11980 21956
rect 12032 21944 12038 21956
rect 14458 21944 14464 21956
rect 12032 21916 14464 21944
rect 12032 21904 12038 21916
rect 14458 21904 14464 21916
rect 14516 21944 14522 21956
rect 14752 21944 14780 21984
rect 14516 21916 14780 21944
rect 15381 21947 15439 21953
rect 14516 21904 14522 21916
rect 15381 21913 15393 21947
rect 15427 21913 15439 21947
rect 15488 21944 15516 21984
rect 15565 21981 15577 22015
rect 15611 22012 15623 22015
rect 16761 22015 16819 22021
rect 16761 22012 16773 22015
rect 15611 21984 16773 22012
rect 15611 21981 15623 21984
rect 15565 21975 15623 21981
rect 16025 21947 16083 21953
rect 16025 21944 16037 21947
rect 15488 21916 16037 21944
rect 15381 21907 15439 21913
rect 16025 21913 16037 21916
rect 16071 21913 16083 21947
rect 16025 21907 16083 21913
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 7708 21848 7849 21876
rect 7708 21836 7714 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 8202 21836 8208 21888
rect 8260 21836 8266 21888
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21876 9551 21879
rect 9674 21876 9680 21888
rect 9539 21848 9680 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10413 21879 10471 21885
rect 10413 21876 10425 21879
rect 9824 21848 10425 21876
rect 9824 21836 9830 21848
rect 10413 21845 10425 21848
rect 10459 21845 10471 21879
rect 10413 21839 10471 21845
rect 11606 21836 11612 21888
rect 11664 21836 11670 21888
rect 11790 21836 11796 21888
rect 11848 21876 11854 21888
rect 15396 21876 15424 21907
rect 11848 21848 15424 21876
rect 11848 21836 11854 21848
rect 15838 21836 15844 21888
rect 15896 21836 15902 21888
rect 16040 21876 16068 21907
rect 16114 21904 16120 21956
rect 16172 21944 16178 21956
rect 16209 21947 16267 21953
rect 16209 21944 16221 21947
rect 16172 21916 16221 21944
rect 16172 21904 16178 21916
rect 16209 21913 16221 21916
rect 16255 21913 16267 21947
rect 16209 21907 16267 21913
rect 16298 21904 16304 21956
rect 16356 21904 16362 21956
rect 16482 21904 16488 21956
rect 16540 21904 16546 21956
rect 16500 21876 16528 21904
rect 16040 21848 16528 21876
rect 16592 21876 16620 21984
rect 16761 21981 16773 21984
rect 16807 21981 16819 22015
rect 16761 21975 16819 21981
rect 16942 21972 16948 22024
rect 17000 21972 17006 22024
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 17313 21975 17371 21981
rect 16669 21947 16727 21953
rect 16669 21913 16681 21947
rect 16715 21944 16727 21947
rect 17319 21944 17347 21975
rect 16715 21916 17347 21944
rect 18984 21944 19012 22188
rect 24394 22108 24400 22160
rect 24452 22108 24458 22160
rect 19245 22083 19303 22089
rect 19245 22049 19257 22083
rect 19291 22080 19303 22083
rect 20530 22080 20536 22092
rect 19291 22052 20536 22080
rect 19291 22049 19303 22052
rect 19245 22043 19303 22049
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 23750 21972 23756 22024
rect 23808 21972 23814 22024
rect 19426 21944 19432 21956
rect 18984 21916 19432 21944
rect 16715 21913 16727 21916
rect 16669 21907 16727 21913
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21944 19579 21947
rect 19794 21944 19800 21956
rect 19567 21916 19800 21944
rect 19567 21913 19579 21916
rect 19521 21907 19579 21913
rect 19794 21904 19800 21916
rect 19852 21904 19858 21956
rect 20162 21904 20168 21956
rect 20220 21904 20226 21956
rect 20824 21916 22094 21944
rect 20824 21876 20852 21916
rect 16592 21848 20852 21876
rect 20990 21836 20996 21888
rect 21048 21836 21054 21888
rect 22066 21876 22094 21916
rect 24026 21904 24032 21956
rect 24084 21944 24090 21956
rect 24302 21944 24308 21956
rect 24084 21916 24308 21944
rect 24084 21904 24090 21916
rect 24302 21904 24308 21916
rect 24360 21904 24366 21956
rect 24581 21947 24639 21953
rect 24581 21913 24593 21947
rect 24627 21913 24639 21947
rect 24581 21907 24639 21913
rect 23937 21879 23995 21885
rect 23937 21876 23949 21879
rect 22066 21848 23949 21876
rect 23937 21845 23949 21848
rect 23983 21876 23995 21879
rect 24596 21876 24624 21907
rect 23983 21848 24624 21876
rect 23983 21845 23995 21848
rect 23937 21839 23995 21845
rect 1104 21786 31280 21808
rect 1104 21734 4922 21786
rect 4974 21734 4986 21786
rect 5038 21734 5050 21786
rect 5102 21734 5114 21786
rect 5166 21734 5178 21786
rect 5230 21734 5242 21786
rect 5294 21734 10922 21786
rect 10974 21734 10986 21786
rect 11038 21734 11050 21786
rect 11102 21734 11114 21786
rect 11166 21734 11178 21786
rect 11230 21734 11242 21786
rect 11294 21734 16922 21786
rect 16974 21734 16986 21786
rect 17038 21734 17050 21786
rect 17102 21734 17114 21786
rect 17166 21734 17178 21786
rect 17230 21734 17242 21786
rect 17294 21734 22922 21786
rect 22974 21734 22986 21786
rect 23038 21734 23050 21786
rect 23102 21734 23114 21786
rect 23166 21734 23178 21786
rect 23230 21734 23242 21786
rect 23294 21734 28922 21786
rect 28974 21734 28986 21786
rect 29038 21734 29050 21786
rect 29102 21734 29114 21786
rect 29166 21734 29178 21786
rect 29230 21734 29242 21786
rect 29294 21734 31280 21786
rect 1104 21712 31280 21734
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 8849 21675 8907 21681
rect 8849 21672 8861 21675
rect 8260 21644 8861 21672
rect 8260 21632 8266 21644
rect 8849 21641 8861 21644
rect 8895 21641 8907 21675
rect 8849 21635 8907 21641
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10100 21644 12434 21672
rect 10100 21632 10106 21644
rect 6549 21607 6607 21613
rect 6549 21573 6561 21607
rect 6595 21604 6607 21607
rect 7374 21604 7380 21616
rect 6595 21576 7380 21604
rect 6595 21573 6607 21576
rect 6549 21567 6607 21573
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 8757 21607 8815 21613
rect 8757 21573 8769 21607
rect 8803 21604 8815 21607
rect 12406 21604 12434 21644
rect 13078 21632 13084 21684
rect 13136 21632 13142 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 14090 21672 14096 21684
rect 13587 21644 14096 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 14090 21632 14096 21644
rect 14148 21632 14154 21684
rect 15838 21632 15844 21684
rect 15896 21632 15902 21684
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 20346 21672 20352 21684
rect 17460 21644 20352 21672
rect 17460 21632 17466 21644
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 15194 21604 15200 21616
rect 8803 21576 10732 21604
rect 12406 21576 15200 21604
rect 8803 21573 8815 21576
rect 8757 21567 8815 21573
rect 10704 21548 10732 21576
rect 15194 21564 15200 21576
rect 15252 21604 15258 21616
rect 15289 21607 15347 21613
rect 15289 21604 15301 21607
rect 15252 21576 15301 21604
rect 15252 21564 15258 21576
rect 15289 21573 15301 21576
rect 15335 21573 15347 21607
rect 15289 21567 15347 21573
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 5997 21471 6055 21477
rect 5997 21468 6009 21471
rect 5184 21440 6009 21468
rect 5184 21344 5212 21440
rect 5997 21437 6009 21440
rect 6043 21468 6055 21471
rect 6380 21468 6408 21499
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 7558 21536 7564 21548
rect 6779 21508 7564 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 9585 21539 9643 21545
rect 9585 21536 9597 21539
rect 8772 21508 9597 21536
rect 8772 21480 8800 21508
rect 9585 21505 9597 21508
rect 9631 21505 9643 21539
rect 9585 21499 9643 21505
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 9841 21539 9899 21545
rect 9841 21536 9853 21539
rect 9732 21508 9853 21536
rect 9732 21496 9738 21508
rect 9841 21505 9853 21508
rect 9887 21505 9899 21539
rect 9841 21499 9899 21505
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 11968 21539 12026 21545
rect 11968 21505 11980 21539
rect 12014 21536 12026 21539
rect 12526 21536 12532 21548
rect 12014 21508 12532 21536
rect 12014 21505 12026 21508
rect 11968 21499 12026 21505
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 15856 21536 15884 21632
rect 16853 21607 16911 21613
rect 16853 21573 16865 21607
rect 16899 21604 16911 21607
rect 16942 21604 16948 21616
rect 16899 21576 16948 21604
rect 16899 21573 16911 21576
rect 16853 21567 16911 21573
rect 16942 21564 16948 21576
rect 17000 21564 17006 21616
rect 17037 21607 17095 21613
rect 17037 21573 17049 21607
rect 17083 21604 17095 21607
rect 18046 21604 18052 21616
rect 17083 21576 18052 21604
rect 17083 21573 17095 21576
rect 17037 21567 17095 21573
rect 18046 21564 18052 21576
rect 18104 21564 18110 21616
rect 21818 21564 21824 21616
rect 21876 21564 21882 21616
rect 15933 21539 15991 21545
rect 15933 21536 15945 21539
rect 15856 21508 15945 21536
rect 15933 21505 15945 21508
rect 15979 21505 15991 21539
rect 15933 21499 15991 21505
rect 16298 21496 16304 21548
rect 16356 21536 16362 21548
rect 17126 21536 17132 21548
rect 16356 21508 17132 21536
rect 16356 21496 16362 21508
rect 17126 21496 17132 21508
rect 17184 21536 17190 21548
rect 17313 21539 17371 21545
rect 17313 21536 17325 21539
rect 17184 21508 17325 21536
rect 17184 21496 17190 21508
rect 17313 21505 17325 21508
rect 17359 21505 17371 21539
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17313 21499 17371 21505
rect 17665 21505 17693 21536
rect 17727 21505 17739 21539
rect 17665 21499 17739 21505
rect 6043 21440 6408 21468
rect 6043 21437 6055 21440
rect 5997 21431 6055 21437
rect 7098 21428 7104 21480
rect 7156 21468 7162 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7156 21440 7941 21468
rect 7156 21428 7162 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 8754 21428 8760 21480
rect 8812 21428 8818 21480
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21437 9551 21471
rect 9493 21431 9551 21437
rect 5166 21292 5172 21344
rect 5224 21292 5230 21344
rect 5442 21292 5448 21344
rect 5500 21292 5506 21344
rect 6917 21335 6975 21341
rect 6917 21301 6929 21335
rect 6963 21332 6975 21335
rect 8294 21332 8300 21344
rect 6963 21304 8300 21332
rect 6963 21301 6975 21304
rect 6917 21295 6975 21301
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 9508 21332 9536 21431
rect 11054 21428 11060 21480
rect 11112 21468 11118 21480
rect 11698 21468 11704 21480
rect 11112 21440 11704 21468
rect 11112 21428 11118 21440
rect 11698 21428 11704 21440
rect 11756 21428 11762 21480
rect 12986 21428 12992 21480
rect 13044 21428 13050 21480
rect 13630 21428 13636 21480
rect 13688 21428 13694 21480
rect 13817 21471 13875 21477
rect 13817 21437 13829 21471
rect 13863 21468 13875 21471
rect 14550 21468 14556 21480
rect 13863 21440 14556 21468
rect 13863 21437 13875 21440
rect 13817 21431 13875 21437
rect 14550 21428 14556 21440
rect 14608 21428 14614 21480
rect 15838 21428 15844 21480
rect 15896 21428 15902 21480
rect 16482 21428 16488 21480
rect 16540 21428 16546 21480
rect 17218 21428 17224 21480
rect 17276 21468 17282 21480
rect 17451 21471 17509 21477
rect 17451 21468 17463 21471
rect 17276 21440 17463 21468
rect 17276 21428 17282 21440
rect 17451 21437 17463 21440
rect 17497 21437 17509 21471
rect 17451 21431 17509 21437
rect 13004 21400 13032 21428
rect 16669 21403 16727 21409
rect 13004 21372 16620 21400
rect 9950 21332 9956 21344
rect 8444 21304 9956 21332
rect 8444 21292 8450 21304
rect 9950 21292 9956 21304
rect 10008 21292 10014 21344
rect 10965 21335 11023 21341
rect 10965 21301 10977 21335
rect 11011 21332 11023 21335
rect 11606 21332 11612 21344
rect 11011 21304 11612 21332
rect 11011 21301 11023 21304
rect 10965 21295 11023 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 13170 21292 13176 21344
rect 13228 21292 13234 21344
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 16482 21332 16488 21344
rect 14792 21304 16488 21332
rect 14792 21292 14798 21304
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 16592 21332 16620 21372
rect 16669 21369 16681 21403
rect 16715 21400 16727 21403
rect 17665 21400 17693 21499
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 21836 21536 21864 21564
rect 17920 21508 21864 21536
rect 17920 21496 17926 21508
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 22152 21508 22201 21536
rect 22152 21496 22158 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 23382 21496 23388 21548
rect 23440 21496 23446 21548
rect 23753 21539 23811 21545
rect 23753 21505 23765 21539
rect 23799 21536 23811 21539
rect 23799 21508 24164 21536
rect 23799 21505 23811 21508
rect 23753 21499 23811 21505
rect 17770 21428 17776 21480
rect 17828 21428 17834 21480
rect 18049 21471 18107 21477
rect 18049 21437 18061 21471
rect 18095 21468 18107 21471
rect 20898 21468 20904 21480
rect 18095 21440 20904 21468
rect 18095 21437 18107 21440
rect 18049 21431 18107 21437
rect 16715 21372 17693 21400
rect 16715 21369 16727 21372
rect 16669 21363 16727 21369
rect 18064 21332 18092 21431
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 23474 21428 23480 21480
rect 23532 21468 23538 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 23532 21440 23673 21468
rect 23532 21428 23538 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23870 21471 23928 21477
rect 23870 21437 23882 21471
rect 23916 21468 23928 21471
rect 24026 21468 24032 21480
rect 23916 21440 24032 21468
rect 23916 21437 23928 21440
rect 23870 21431 23928 21437
rect 24026 21428 24032 21440
rect 24084 21428 24090 21480
rect 24136 21400 24164 21508
rect 24210 21496 24216 21548
rect 24268 21496 24274 21548
rect 24136 21372 24440 21400
rect 24412 21344 24440 21372
rect 16592 21304 18092 21332
rect 24029 21335 24087 21341
rect 24029 21301 24041 21335
rect 24075 21332 24087 21335
rect 24210 21332 24216 21344
rect 24075 21304 24216 21332
rect 24075 21301 24087 21304
rect 24029 21295 24087 21301
rect 24210 21292 24216 21304
rect 24268 21292 24274 21344
rect 24302 21292 24308 21344
rect 24360 21292 24366 21344
rect 24394 21292 24400 21344
rect 24452 21292 24458 21344
rect 1104 21242 31280 21264
rect 1104 21190 4182 21242
rect 4234 21190 4246 21242
rect 4298 21190 4310 21242
rect 4362 21190 4374 21242
rect 4426 21190 4438 21242
rect 4490 21190 4502 21242
rect 4554 21190 10182 21242
rect 10234 21190 10246 21242
rect 10298 21190 10310 21242
rect 10362 21190 10374 21242
rect 10426 21190 10438 21242
rect 10490 21190 10502 21242
rect 10554 21190 16182 21242
rect 16234 21190 16246 21242
rect 16298 21190 16310 21242
rect 16362 21190 16374 21242
rect 16426 21190 16438 21242
rect 16490 21190 16502 21242
rect 16554 21190 22182 21242
rect 22234 21190 22246 21242
rect 22298 21190 22310 21242
rect 22362 21190 22374 21242
rect 22426 21190 22438 21242
rect 22490 21190 22502 21242
rect 22554 21190 28182 21242
rect 28234 21190 28246 21242
rect 28298 21190 28310 21242
rect 28362 21190 28374 21242
rect 28426 21190 28438 21242
rect 28490 21190 28502 21242
rect 28554 21190 31280 21242
rect 1104 21168 31280 21190
rect 5166 21088 5172 21140
rect 5224 21088 5230 21140
rect 5442 21088 5448 21140
rect 5500 21128 5506 21140
rect 5500 21100 5672 21128
rect 5500 21088 5506 21100
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20924 3847 20927
rect 3878 20924 3884 20936
rect 3835 20896 3884 20924
rect 3835 20893 3847 20896
rect 3789 20887 3847 20893
rect 3878 20884 3884 20896
rect 3936 20924 3942 20936
rect 5644 20933 5672 21100
rect 6288 21100 7972 21128
rect 5902 20952 5908 21004
rect 5960 20992 5966 21004
rect 6288 20992 6316 21100
rect 7944 21060 7972 21100
rect 8386 21088 8392 21140
rect 8444 21088 8450 21140
rect 9306 21088 9312 21140
rect 9364 21128 9370 21140
rect 9401 21131 9459 21137
rect 9401 21128 9413 21131
rect 9364 21100 9413 21128
rect 9364 21088 9370 21100
rect 9401 21097 9413 21100
rect 9447 21097 9459 21131
rect 9401 21091 9459 21097
rect 12526 21088 12532 21140
rect 12584 21088 12590 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13170 21088 13176 21140
rect 13228 21088 13234 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 17218 21128 17224 21140
rect 13320 21100 17224 21128
rect 13320 21088 13326 21100
rect 17218 21088 17224 21100
rect 17276 21128 17282 21140
rect 17862 21128 17868 21140
rect 17276 21100 17868 21128
rect 17276 21088 17282 21100
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19521 21131 19579 21137
rect 19521 21128 19533 21131
rect 19392 21100 19533 21128
rect 19392 21088 19398 21100
rect 19521 21097 19533 21100
rect 19567 21128 19579 21131
rect 19978 21128 19984 21140
rect 19567 21100 19984 21128
rect 19567 21097 19579 21100
rect 19521 21091 19579 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 20162 21088 20168 21140
rect 20220 21088 20226 21140
rect 22094 21088 22100 21140
rect 22152 21128 22158 21140
rect 22373 21131 22431 21137
rect 22373 21128 22385 21131
rect 22152 21100 22385 21128
rect 22152 21088 22158 21100
rect 22373 21097 22385 21100
rect 22419 21097 22431 21131
rect 22373 21091 22431 21097
rect 23661 21131 23719 21137
rect 23661 21097 23673 21131
rect 23707 21128 23719 21131
rect 23750 21128 23756 21140
rect 23707 21100 23756 21128
rect 23707 21097 23719 21100
rect 23661 21091 23719 21097
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 23934 21088 23940 21140
rect 23992 21128 23998 21140
rect 24489 21131 24547 21137
rect 24489 21128 24501 21131
rect 23992 21100 24501 21128
rect 23992 21088 23998 21100
rect 24489 21097 24501 21100
rect 24535 21097 24547 21131
rect 24489 21091 24547 21097
rect 12986 21060 12992 21072
rect 7944 21032 12992 21060
rect 12986 21020 12992 21032
rect 13044 21020 13050 21072
rect 5960 20964 6316 20992
rect 6365 20995 6423 21001
rect 5960 20952 5966 20964
rect 6365 20961 6377 20995
rect 6411 20992 6423 20995
rect 6638 20992 6644 21004
rect 6411 20964 6644 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 8110 20952 8116 21004
rect 8168 20992 8174 21004
rect 9861 20995 9919 21001
rect 9861 20992 9873 20995
rect 8168 20964 9873 20992
rect 8168 20952 8174 20964
rect 9861 20961 9873 20964
rect 9907 20961 9919 20995
rect 9861 20955 9919 20961
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 13096 20992 13124 21088
rect 11900 20964 13124 20992
rect 5629 20927 5687 20933
rect 3936 20896 4844 20924
rect 3936 20884 3942 20896
rect 4816 20868 4844 20896
rect 5629 20893 5641 20927
rect 5675 20893 5687 20927
rect 5629 20887 5687 20893
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20924 7067 20927
rect 7098 20924 7104 20936
rect 7055 20896 7104 20924
rect 7055 20893 7067 20896
rect 7009 20887 7067 20893
rect 4056 20859 4114 20865
rect 4056 20825 4068 20859
rect 4102 20856 4114 20859
rect 4154 20856 4160 20868
rect 4102 20828 4160 20856
rect 4102 20825 4114 20828
rect 4056 20819 4114 20825
rect 4154 20816 4160 20828
rect 4212 20816 4218 20868
rect 4798 20816 4804 20868
rect 4856 20856 4862 20868
rect 7024 20856 7052 20887
rect 7098 20884 7104 20896
rect 7156 20884 7162 20936
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 9674 20924 9680 20936
rect 8803 20896 9680 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 9674 20884 9680 20896
rect 9732 20884 9738 20936
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 10229 20927 10287 20933
rect 10229 20893 10241 20927
rect 10275 20924 10287 20927
rect 10686 20924 10692 20936
rect 10275 20896 10692 20924
rect 10275 20893 10287 20896
rect 10229 20887 10287 20893
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 11422 20884 11428 20936
rect 11480 20884 11486 20936
rect 11606 20884 11612 20936
rect 11664 20884 11670 20936
rect 11900 20933 11928 20964
rect 11885 20927 11943 20933
rect 11885 20893 11897 20927
rect 11931 20893 11943 20927
rect 11885 20887 11943 20893
rect 11974 20884 11980 20936
rect 12032 20884 12038 20936
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 12618 20924 12624 20936
rect 12483 20896 12624 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20924 12771 20927
rect 13188 20924 13216 21088
rect 15838 21020 15844 21072
rect 15896 21060 15902 21072
rect 24302 21060 24308 21072
rect 15896 21032 16712 21060
rect 15896 21020 15902 21032
rect 13722 20952 13728 21004
rect 13780 20992 13786 21004
rect 16132 21001 16160 21032
rect 16684 21004 16712 21032
rect 17328 21032 18000 21060
rect 15381 20995 15439 21001
rect 15381 20992 15393 20995
rect 13780 20964 15393 20992
rect 13780 20952 13786 20964
rect 15381 20961 15393 20964
rect 15427 20961 15439 20995
rect 15381 20955 15439 20961
rect 16117 20995 16175 21001
rect 16117 20961 16129 20995
rect 16163 20961 16175 20995
rect 16117 20955 16175 20961
rect 16224 20964 16528 20992
rect 12759 20896 13216 20924
rect 12759 20893 12771 20896
rect 12713 20887 12771 20893
rect 14642 20884 14648 20936
rect 14700 20884 14706 20936
rect 16022 20884 16028 20936
rect 16080 20884 16086 20936
rect 4856 20828 7052 20856
rect 7276 20859 7334 20865
rect 4856 20816 4862 20828
rect 7276 20825 7288 20859
rect 7322 20856 7334 20859
rect 7466 20856 7472 20868
rect 7322 20828 7472 20856
rect 7322 20825 7334 20828
rect 7276 20819 7334 20825
rect 7466 20816 7472 20828
rect 7524 20816 7530 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 8772 20828 10977 20856
rect 8772 20800 8800 20828
rect 10965 20825 10977 20828
rect 11011 20856 11023 20859
rect 11054 20856 11060 20868
rect 11011 20828 11060 20856
rect 11011 20825 11023 20828
rect 10965 20819 11023 20825
rect 11054 20816 11060 20828
rect 11112 20816 11118 20868
rect 11440 20856 11468 20884
rect 11793 20859 11851 20865
rect 11793 20856 11805 20859
rect 11440 20828 11805 20856
rect 11793 20825 11805 20828
rect 11839 20825 11851 20859
rect 11793 20819 11851 20825
rect 15286 20816 15292 20868
rect 15344 20856 15350 20868
rect 16224 20856 16252 20964
rect 16500 20936 16528 20964
rect 16666 20952 16672 21004
rect 16724 20952 16730 21004
rect 16758 20952 16764 21004
rect 16816 20952 16822 21004
rect 16942 20952 16948 21004
rect 17000 20992 17006 21004
rect 17328 20992 17356 21032
rect 17000 20964 17356 20992
rect 17405 20995 17463 21001
rect 17000 20952 17006 20964
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17494 20992 17500 21004
rect 17451 20964 17500 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 17865 20995 17923 21001
rect 17865 20961 17877 20995
rect 17911 20992 17923 20995
rect 17972 20992 18000 21032
rect 19306 21032 24308 21060
rect 19306 20992 19334 21032
rect 24302 21020 24308 21032
rect 24360 21020 24366 21072
rect 17911 20964 19334 20992
rect 17911 20961 17923 20964
rect 17865 20955 17923 20961
rect 19610 20952 19616 21004
rect 19668 20992 19674 21004
rect 20717 20995 20775 21001
rect 20717 20992 20729 20995
rect 19668 20964 20729 20992
rect 19668 20952 19674 20964
rect 20717 20961 20729 20964
rect 20763 20961 20775 20995
rect 22214 20995 22272 21001
rect 22214 20992 22226 20995
rect 20717 20955 20775 20961
rect 21100 20964 22226 20992
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 15344 20828 16252 20856
rect 16408 20856 16436 20887
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16577 20927 16635 20933
rect 16577 20924 16589 20927
rect 16540 20896 16589 20924
rect 16540 20884 16546 20896
rect 16577 20893 16589 20896
rect 16623 20893 16635 20927
rect 16577 20887 16635 20893
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17328 20856 17356 20887
rect 17678 20884 17684 20936
rect 17736 20884 17742 20936
rect 18046 20884 18052 20936
rect 18104 20924 18110 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18104 20896 18429 20924
rect 18104 20884 18110 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20924 20683 20927
rect 20990 20924 20996 20936
rect 20671 20896 20996 20924
rect 20671 20893 20683 20896
rect 20625 20887 20683 20893
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21100 20933 21128 20964
rect 22214 20961 22226 20964
rect 22260 20992 22272 20995
rect 22462 20992 22468 21004
rect 22260 20964 22468 20992
rect 22260 20961 22272 20964
rect 22214 20955 22272 20961
rect 22462 20952 22468 20964
rect 22520 20952 22526 21004
rect 23382 20952 23388 21004
rect 23440 20952 23446 21004
rect 23474 20952 23480 21004
rect 23532 20992 23538 21004
rect 23532 20964 23888 20992
rect 23532 20952 23538 20964
rect 21085 20927 21143 20933
rect 21085 20893 21097 20927
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 21634 20884 21640 20936
rect 21692 20884 21698 20936
rect 21726 20884 21732 20936
rect 21784 20884 21790 20936
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21928 20896 22017 20924
rect 17957 20859 18015 20865
rect 17957 20856 17969 20859
rect 16408 20828 17172 20856
rect 17328 20828 17969 20856
rect 15344 20816 15350 20828
rect 17144 20800 17172 20828
rect 17957 20825 17969 20828
rect 18003 20825 18015 20859
rect 17957 20819 18015 20825
rect 18141 20859 18199 20865
rect 18141 20825 18153 20859
rect 18187 20856 18199 20859
rect 18230 20856 18236 20868
rect 18187 20828 18236 20856
rect 18187 20825 18199 20828
rect 18141 20819 18199 20825
rect 18230 20816 18236 20828
rect 18288 20816 18294 20868
rect 18322 20816 18328 20868
rect 18380 20856 18386 20868
rect 18380 20828 18644 20856
rect 18380 20816 18386 20828
rect 5261 20791 5319 20797
rect 5261 20757 5273 20791
rect 5307 20788 5319 20791
rect 5350 20788 5356 20800
rect 5307 20760 5356 20788
rect 5307 20757 5319 20760
rect 5261 20751 5319 20757
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 5718 20748 5724 20800
rect 5776 20748 5782 20800
rect 6914 20748 6920 20800
rect 6972 20748 6978 20800
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8573 20791 8631 20797
rect 8573 20788 8585 20791
rect 8536 20760 8585 20788
rect 8536 20748 8542 20760
rect 8573 20757 8585 20760
rect 8619 20757 8631 20791
rect 8573 20751 8631 20757
rect 8754 20748 8760 20800
rect 8812 20748 8818 20800
rect 11422 20748 11428 20800
rect 11480 20788 11486 20800
rect 12161 20791 12219 20797
rect 12161 20788 12173 20791
rect 11480 20760 12173 20788
rect 11480 20748 11486 20760
rect 12161 20757 12173 20760
rect 12207 20757 12219 20791
rect 12161 20751 12219 20757
rect 12250 20748 12256 20800
rect 12308 20748 12314 20800
rect 14090 20748 14096 20800
rect 14148 20748 14154 20800
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17678 20788 17684 20800
rect 17184 20760 17684 20788
rect 17184 20748 17190 20760
rect 17678 20748 17684 20760
rect 17736 20748 17742 20800
rect 18616 20797 18644 20828
rect 19058 20816 19064 20868
rect 19116 20856 19122 20868
rect 19429 20859 19487 20865
rect 19429 20856 19441 20859
rect 19116 20828 19441 20856
rect 19116 20816 19122 20828
rect 19429 20825 19441 20828
rect 19475 20825 19487 20859
rect 19429 20819 19487 20825
rect 21177 20859 21235 20865
rect 21177 20825 21189 20859
rect 21223 20856 21235 20859
rect 21928 20856 21956 20896
rect 22005 20893 22017 20896
rect 22051 20924 22063 20927
rect 23017 20927 23075 20933
rect 23017 20924 23029 20927
rect 22051 20896 23029 20924
rect 22051 20893 22063 20896
rect 22005 20887 22063 20893
rect 23017 20893 23029 20896
rect 23063 20924 23075 20927
rect 23400 20924 23428 20952
rect 23750 20924 23756 20936
rect 23063 20896 23756 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 23750 20884 23756 20896
rect 23808 20884 23814 20936
rect 23860 20933 23888 20964
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20893 23903 20927
rect 23845 20887 23903 20893
rect 23934 20884 23940 20936
rect 23992 20884 23998 20936
rect 24026 20884 24032 20936
rect 24084 20884 24090 20936
rect 24121 20927 24179 20933
rect 24121 20893 24133 20927
rect 24167 20924 24179 20927
rect 24394 20924 24400 20936
rect 24167 20896 24400 20924
rect 24167 20893 24179 20896
rect 24121 20887 24179 20893
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 21223 20828 21956 20856
rect 21223 20825 21235 20828
rect 21177 20819 21235 20825
rect 23382 20816 23388 20868
rect 23440 20856 23446 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 23440 20828 24593 20856
rect 23440 20816 23446 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24581 20819 24639 20825
rect 18601 20791 18659 20797
rect 18601 20757 18613 20791
rect 18647 20757 18659 20791
rect 18601 20751 18659 20757
rect 21634 20748 21640 20800
rect 21692 20788 21698 20800
rect 22097 20791 22155 20797
rect 22097 20788 22109 20791
rect 21692 20760 22109 20788
rect 21692 20748 21698 20760
rect 22097 20757 22109 20760
rect 22143 20757 22155 20791
rect 22097 20751 22155 20757
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 22554 20788 22560 20800
rect 22244 20760 22560 20788
rect 22244 20748 22250 20760
rect 22554 20748 22560 20760
rect 22612 20788 22618 20800
rect 22925 20791 22983 20797
rect 22925 20788 22937 20791
rect 22612 20760 22937 20788
rect 22612 20748 22618 20760
rect 22925 20757 22937 20760
rect 22971 20788 22983 20791
rect 23658 20788 23664 20800
rect 22971 20760 23664 20788
rect 22971 20757 22983 20760
rect 22925 20751 22983 20757
rect 23658 20748 23664 20760
rect 23716 20788 23722 20800
rect 23934 20788 23940 20800
rect 23716 20760 23940 20788
rect 23716 20748 23722 20760
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 1104 20698 31280 20720
rect 1104 20646 4922 20698
rect 4974 20646 4986 20698
rect 5038 20646 5050 20698
rect 5102 20646 5114 20698
rect 5166 20646 5178 20698
rect 5230 20646 5242 20698
rect 5294 20646 10922 20698
rect 10974 20646 10986 20698
rect 11038 20646 11050 20698
rect 11102 20646 11114 20698
rect 11166 20646 11178 20698
rect 11230 20646 11242 20698
rect 11294 20646 16922 20698
rect 16974 20646 16986 20698
rect 17038 20646 17050 20698
rect 17102 20646 17114 20698
rect 17166 20646 17178 20698
rect 17230 20646 17242 20698
rect 17294 20646 22922 20698
rect 22974 20646 22986 20698
rect 23038 20646 23050 20698
rect 23102 20646 23114 20698
rect 23166 20646 23178 20698
rect 23230 20646 23242 20698
rect 23294 20646 28922 20698
rect 28974 20646 28986 20698
rect 29038 20646 29050 20698
rect 29102 20646 29114 20698
rect 29166 20646 29178 20698
rect 29230 20646 29242 20698
rect 29294 20646 31280 20698
rect 1104 20624 31280 20646
rect 4154 20544 4160 20596
rect 4212 20544 4218 20596
rect 5350 20544 5356 20596
rect 5408 20544 5414 20596
rect 6181 20587 6239 20593
rect 6181 20553 6193 20587
rect 6227 20584 6239 20587
rect 6638 20584 6644 20596
rect 6227 20556 6644 20584
rect 6227 20553 6239 20556
rect 6181 20547 6239 20553
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 6825 20587 6883 20593
rect 6825 20553 6837 20587
rect 6871 20584 6883 20587
rect 6914 20584 6920 20596
rect 6871 20556 6920 20584
rect 6871 20553 6883 20556
rect 6825 20547 6883 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 7466 20544 7472 20596
rect 7524 20544 7530 20596
rect 9585 20587 9643 20593
rect 8128 20556 8892 20584
rect 5368 20516 5396 20544
rect 8128 20516 8156 20556
rect 4356 20488 5396 20516
rect 6748 20488 8156 20516
rect 8220 20488 8800 20516
rect 4356 20457 4384 20488
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 5068 20451 5126 20457
rect 5068 20417 5080 20451
rect 5114 20448 5126 20451
rect 5534 20448 5540 20460
rect 5114 20420 5540 20448
rect 5114 20417 5126 20420
rect 5068 20411 5126 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6748 20457 6776 20488
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6144 20420 6745 20448
rect 6144 20408 6150 20420
rect 6733 20417 6745 20420
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 7650 20408 7656 20460
rect 7708 20408 7714 20460
rect 8220 20457 8248 20488
rect 8772 20460 8800 20488
rect 8478 20457 8484 20460
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8472 20448 8484 20457
rect 8439 20420 8484 20448
rect 8205 20411 8263 20417
rect 8472 20411 8484 20420
rect 8478 20408 8484 20411
rect 8536 20408 8542 20460
rect 8754 20408 8760 20460
rect 8812 20408 8818 20460
rect 8864 20448 8892 20556
rect 9585 20553 9597 20587
rect 9631 20553 9643 20587
rect 9585 20547 9643 20553
rect 9600 20516 9628 20547
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 11164 20556 12572 20584
rect 9600 20488 11100 20516
rect 10796 20460 10824 20488
rect 10045 20451 10103 20457
rect 8864 20420 9260 20448
rect 4798 20340 4804 20392
rect 4856 20340 4862 20392
rect 6822 20340 6828 20392
rect 6880 20380 6886 20392
rect 6917 20383 6975 20389
rect 6917 20380 6929 20383
rect 6880 20352 6929 20380
rect 6880 20340 6886 20352
rect 6917 20349 6929 20352
rect 6963 20349 6975 20383
rect 9232 20380 9260 20420
rect 10045 20417 10057 20451
rect 10091 20448 10103 20451
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10091 20420 10517 20448
rect 10091 20417 10103 20420
rect 10045 20411 10103 20417
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 10778 20408 10784 20460
rect 10836 20408 10842 20460
rect 11072 20457 11100 20488
rect 11057 20451 11115 20457
rect 11057 20417 11069 20451
rect 11103 20417 11115 20451
rect 11057 20411 11115 20417
rect 10137 20383 10195 20389
rect 10137 20380 10149 20383
rect 9232 20352 10149 20380
rect 6917 20343 6975 20349
rect 10137 20349 10149 20352
rect 10183 20349 10195 20383
rect 10137 20343 10195 20349
rect 1854 20272 1860 20324
rect 1912 20272 1918 20324
rect 10152 20312 10180 20343
rect 10318 20340 10324 20392
rect 10376 20340 10382 20392
rect 11164 20312 11192 20556
rect 12434 20516 12440 20528
rect 11900 20488 12440 20516
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 11900 20457 11928 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 12544 20516 12572 20556
rect 12618 20544 12624 20596
rect 12676 20584 12682 20596
rect 13357 20587 13415 20593
rect 13357 20584 13369 20587
rect 12676 20556 13369 20584
rect 12676 20544 12682 20556
rect 13357 20553 13369 20556
rect 13403 20553 13415 20587
rect 13357 20547 13415 20553
rect 13725 20587 13783 20593
rect 13725 20553 13737 20587
rect 13771 20584 13783 20587
rect 14090 20584 14096 20596
rect 13771 20556 14096 20584
rect 13771 20553 13783 20556
rect 13725 20547 13783 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16022 20584 16028 20596
rect 15979 20556 16028 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 18046 20544 18052 20596
rect 18104 20584 18110 20596
rect 18325 20587 18383 20593
rect 18325 20584 18337 20587
rect 18104 20556 18337 20584
rect 18104 20544 18110 20556
rect 14369 20519 14427 20525
rect 12544 20488 13676 20516
rect 12158 20457 12164 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11756 20420 11897 20448
rect 11756 20408 11762 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 12152 20448 12164 20457
rect 12119 20420 12164 20448
rect 11885 20411 11943 20417
rect 12152 20411 12164 20420
rect 12158 20408 12164 20411
rect 12216 20408 12222 20460
rect 13648 20392 13676 20488
rect 14369 20485 14381 20519
rect 14415 20516 14427 20519
rect 16132 20516 16160 20544
rect 16301 20519 16359 20525
rect 16301 20516 16313 20519
rect 14415 20488 14872 20516
rect 14415 20485 14427 20488
rect 14369 20479 14427 20485
rect 14844 20460 14872 20488
rect 15580 20488 16313 20516
rect 15580 20460 15608 20488
rect 16301 20485 16313 20488
rect 16347 20485 16359 20519
rect 16301 20479 16359 20485
rect 16666 20476 16672 20528
rect 16724 20516 16730 20528
rect 17037 20519 17095 20525
rect 17037 20516 17049 20519
rect 16724 20488 17049 20516
rect 16724 20476 16730 20488
rect 17037 20485 17049 20488
rect 17083 20516 17095 20519
rect 17586 20516 17592 20528
rect 17083 20488 17592 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 17586 20476 17592 20488
rect 17644 20476 17650 20528
rect 18248 20525 18276 20556
rect 18325 20553 18337 20556
rect 18371 20553 18383 20587
rect 21542 20584 21548 20596
rect 18325 20547 18383 20553
rect 18432 20556 18736 20584
rect 18233 20519 18291 20525
rect 17696 20488 18184 20516
rect 13722 20408 13728 20460
rect 13780 20448 13786 20460
rect 13780 20420 13952 20448
rect 13780 20408 13786 20420
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 13924 20389 13952 20420
rect 14642 20408 14648 20460
rect 14700 20408 14706 20460
rect 14734 20408 14740 20460
rect 14792 20408 14798 20460
rect 14826 20408 14832 20460
rect 14884 20408 14890 20460
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 15562 20448 15568 20460
rect 15519 20420 15568 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15657 20451 15715 20457
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 13817 20383 13875 20389
rect 13817 20380 13829 20383
rect 13688 20352 13829 20380
rect 13688 20340 13694 20352
rect 13817 20349 13829 20352
rect 13863 20349 13875 20383
rect 13817 20343 13875 20349
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 14182 20340 14188 20392
rect 14240 20340 14246 20392
rect 6288 20284 6500 20312
rect 1872 20244 1900 20272
rect 6288 20244 6316 20284
rect 1872 20216 6316 20244
rect 6362 20204 6368 20256
rect 6420 20204 6426 20256
rect 6472 20244 6500 20284
rect 9140 20284 9720 20312
rect 10152 20284 11192 20312
rect 13265 20315 13323 20321
rect 9140 20244 9168 20284
rect 6472 20216 9168 20244
rect 9692 20244 9720 20284
rect 13265 20281 13277 20315
rect 13311 20312 13323 20315
rect 13998 20312 14004 20324
rect 13311 20284 14004 20312
rect 13311 20281 13323 20284
rect 13265 20275 13323 20281
rect 13998 20272 14004 20284
rect 14056 20312 14062 20324
rect 14660 20312 14688 20408
rect 14752 20380 14780 20408
rect 15672 20380 15700 20411
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 16080 20420 16129 20448
rect 16080 20408 16086 20420
rect 16117 20417 16129 20420
rect 16163 20417 16175 20451
rect 17696 20448 17724 20488
rect 16117 20411 16175 20417
rect 16408 20420 17724 20448
rect 16408 20380 16436 20420
rect 17770 20408 17776 20460
rect 17828 20408 17834 20460
rect 17862 20408 17868 20460
rect 17920 20448 17926 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17920 20420 18061 20448
rect 17920 20408 17926 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18156 20448 18184 20488
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 18279 20488 18313 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 18432 20448 18460 20556
rect 18488 20519 18546 20525
rect 18488 20485 18500 20519
rect 18534 20516 18546 20519
rect 18598 20516 18604 20528
rect 18534 20488 18604 20516
rect 18534 20485 18546 20488
rect 18488 20479 18546 20485
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18708 20525 18736 20556
rect 21192 20556 21548 20584
rect 18693 20519 18751 20525
rect 18693 20485 18705 20519
rect 18739 20516 18751 20519
rect 19242 20516 19248 20528
rect 18739 20488 19248 20516
rect 18739 20485 18751 20488
rect 18693 20479 18751 20485
rect 19242 20476 19248 20488
rect 19300 20476 19306 20528
rect 20714 20476 20720 20528
rect 20772 20476 20778 20528
rect 20990 20476 20996 20528
rect 21048 20516 21054 20528
rect 21192 20525 21220 20556
rect 21542 20544 21548 20556
rect 21600 20584 21606 20596
rect 21726 20584 21732 20596
rect 21600 20556 21732 20584
rect 21600 20544 21606 20556
rect 21726 20544 21732 20556
rect 21784 20544 21790 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22186 20584 22192 20596
rect 21876 20556 22192 20584
rect 21876 20544 21882 20556
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 23290 20544 23296 20596
rect 23348 20584 23354 20596
rect 24118 20584 24124 20596
rect 23348 20556 24124 20584
rect 23348 20544 23354 20556
rect 24118 20544 24124 20556
rect 24176 20544 24182 20596
rect 24949 20587 25007 20593
rect 24949 20553 24961 20587
rect 24995 20584 25007 20587
rect 24995 20556 25176 20584
rect 24995 20553 25007 20556
rect 24949 20547 25007 20553
rect 21177 20519 21235 20525
rect 21177 20516 21189 20519
rect 21048 20488 21189 20516
rect 21048 20476 21054 20488
rect 21177 20485 21189 20488
rect 21223 20485 21235 20519
rect 21177 20479 21235 20485
rect 21744 20488 23704 20516
rect 18156 20420 18460 20448
rect 20625 20451 20683 20457
rect 18049 20411 18107 20417
rect 20625 20417 20637 20451
rect 20671 20448 20683 20451
rect 21085 20451 21143 20457
rect 20671 20420 20944 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 20916 20392 20944 20420
rect 21085 20417 21097 20451
rect 21131 20448 21143 20451
rect 21358 20448 21364 20460
rect 21131 20420 21364 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 21744 20392 21772 20488
rect 21910 20448 21916 20460
rect 21836 20420 21916 20448
rect 14752 20352 15700 20380
rect 15948 20352 16436 20380
rect 15948 20312 15976 20352
rect 16482 20340 16488 20392
rect 16540 20380 16546 20392
rect 16540 20352 20760 20380
rect 16540 20340 16546 20352
rect 14056 20284 14688 20312
rect 15764 20284 15976 20312
rect 16040 20284 18552 20312
rect 14056 20272 14062 20284
rect 15764 20244 15792 20284
rect 16040 20256 16068 20284
rect 9692 20216 15792 20244
rect 15838 20204 15844 20256
rect 15896 20204 15902 20256
rect 16022 20204 16028 20256
rect 16080 20204 16086 20256
rect 17494 20204 17500 20256
rect 17552 20244 17558 20256
rect 17770 20244 17776 20256
rect 17552 20216 17776 20244
rect 17552 20204 17558 20216
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 17862 20204 17868 20256
rect 17920 20204 17926 20256
rect 18524 20253 18552 20284
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 19702 20244 19708 20256
rect 18555 20216 19708 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 19702 20204 19708 20216
rect 19760 20204 19766 20256
rect 20732 20244 20760 20352
rect 20898 20340 20904 20392
rect 20956 20340 20962 20392
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20380 21695 20383
rect 21726 20380 21732 20392
rect 21683 20352 21732 20380
rect 21683 20349 21695 20352
rect 21637 20343 21695 20349
rect 21726 20340 21732 20352
rect 21784 20340 21790 20392
rect 20806 20272 20812 20324
rect 20864 20312 20870 20324
rect 21836 20312 21864 20420
rect 21910 20408 21916 20420
rect 21968 20448 21974 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22373 20451 22431 20457
rect 22373 20417 22385 20451
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 22152 20352 22293 20380
rect 22152 20340 22158 20352
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 22388 20380 22416 20411
rect 22554 20408 22560 20460
rect 22612 20408 22618 20460
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20448 23075 20451
rect 23474 20448 23480 20460
rect 23063 20420 23480 20448
rect 23063 20417 23075 20420
rect 23017 20411 23075 20417
rect 23474 20408 23480 20420
rect 23532 20408 23538 20460
rect 23676 20457 23704 20488
rect 23750 20476 23756 20528
rect 23808 20516 23814 20528
rect 25148 20525 25176 20556
rect 25133 20519 25191 20525
rect 23808 20488 24716 20516
rect 23808 20476 23814 20488
rect 24688 20460 24716 20488
rect 25133 20485 25145 20519
rect 25179 20485 25191 20519
rect 25133 20479 25191 20485
rect 23661 20451 23719 20457
rect 23661 20417 23673 20451
rect 23707 20448 23719 20451
rect 24026 20448 24032 20460
rect 23707 20420 24032 20448
rect 23707 20417 23719 20420
rect 23661 20411 23719 20417
rect 24026 20408 24032 20420
rect 24084 20448 24090 20460
rect 24581 20451 24639 20457
rect 24581 20448 24593 20451
rect 24084 20420 24593 20448
rect 24084 20408 24090 20420
rect 24581 20417 24593 20420
rect 24627 20417 24639 20451
rect 24581 20411 24639 20417
rect 24670 20408 24676 20460
rect 24728 20408 24734 20460
rect 23106 20380 23112 20392
rect 22388 20352 23112 20380
rect 22281 20343 22339 20349
rect 23106 20340 23112 20352
rect 23164 20380 23170 20392
rect 23201 20383 23259 20389
rect 23201 20380 23213 20383
rect 23164 20352 23213 20380
rect 23164 20340 23170 20352
rect 23201 20349 23213 20352
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 23290 20340 23296 20392
rect 23348 20340 23354 20392
rect 23492 20380 23520 20408
rect 24213 20383 24271 20389
rect 24213 20380 24225 20383
rect 23492 20352 24225 20380
rect 24213 20349 24225 20352
rect 24259 20349 24271 20383
rect 24213 20343 24271 20349
rect 24305 20383 24363 20389
rect 24305 20349 24317 20383
rect 24351 20380 24363 20383
rect 24394 20380 24400 20392
rect 24351 20352 24400 20380
rect 24351 20349 24363 20352
rect 24305 20343 24363 20349
rect 24394 20340 24400 20352
rect 24452 20340 24458 20392
rect 24790 20383 24848 20389
rect 24790 20380 24802 20383
rect 24668 20352 24802 20380
rect 23308 20312 23336 20340
rect 20864 20284 21864 20312
rect 22388 20284 23336 20312
rect 20864 20272 20870 20284
rect 22388 20244 22416 20284
rect 23566 20272 23572 20324
rect 23624 20312 23630 20324
rect 24668 20312 24696 20352
rect 24790 20349 24802 20352
rect 24836 20349 24848 20383
rect 24790 20343 24848 20349
rect 23624 20284 24696 20312
rect 23624 20272 23630 20284
rect 20732 20216 22416 20244
rect 22462 20204 22468 20256
rect 22520 20244 22526 20256
rect 22922 20244 22928 20256
rect 22520 20216 22928 20244
rect 22520 20204 22526 20216
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 25225 20247 25283 20253
rect 25225 20244 25237 20247
rect 23808 20216 25237 20244
rect 23808 20204 23814 20216
rect 25225 20213 25237 20216
rect 25271 20213 25283 20247
rect 25225 20207 25283 20213
rect 1104 20154 31280 20176
rect 1104 20102 4182 20154
rect 4234 20102 4246 20154
rect 4298 20102 4310 20154
rect 4362 20102 4374 20154
rect 4426 20102 4438 20154
rect 4490 20102 4502 20154
rect 4554 20102 10182 20154
rect 10234 20102 10246 20154
rect 10298 20102 10310 20154
rect 10362 20102 10374 20154
rect 10426 20102 10438 20154
rect 10490 20102 10502 20154
rect 10554 20102 16182 20154
rect 16234 20102 16246 20154
rect 16298 20102 16310 20154
rect 16362 20102 16374 20154
rect 16426 20102 16438 20154
rect 16490 20102 16502 20154
rect 16554 20102 22182 20154
rect 22234 20102 22246 20154
rect 22298 20102 22310 20154
rect 22362 20102 22374 20154
rect 22426 20102 22438 20154
rect 22490 20102 22502 20154
rect 22554 20102 28182 20154
rect 28234 20102 28246 20154
rect 28298 20102 28310 20154
rect 28362 20102 28374 20154
rect 28426 20102 28438 20154
rect 28490 20102 28502 20154
rect 28554 20102 31280 20154
rect 1104 20080 31280 20102
rect 5534 20000 5540 20052
rect 5592 20000 5598 20052
rect 6362 20000 6368 20052
rect 6420 20000 6426 20052
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 6880 20012 11192 20040
rect 6880 20000 6886 20012
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 6380 19836 6408 20000
rect 10778 19932 10784 19984
rect 10836 19932 10842 19984
rect 11057 19975 11115 19981
rect 11057 19941 11069 19975
rect 11103 19941 11115 19975
rect 11164 19972 11192 20012
rect 11422 20000 11428 20052
rect 11480 20000 11486 20052
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 16666 20040 16672 20052
rect 12768 20012 16672 20040
rect 12768 20000 12774 20012
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 18923 20012 19257 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 22094 20040 22100 20052
rect 19245 20003 19303 20009
rect 19536 20012 22100 20040
rect 11164 19944 15700 19972
rect 11057 19935 11115 19941
rect 5767 19808 6408 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 8294 19796 8300 19848
rect 8352 19796 8358 19848
rect 9950 19796 9956 19848
rect 10008 19836 10014 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 10008 19808 10517 19836
rect 10008 19796 10014 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 10796 19845 10824 19932
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10652 19808 10701 19836
rect 10652 19796 10658 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10870 19796 10876 19848
rect 10928 19796 10934 19848
rect 11072 19836 11100 19935
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 11379 19876 12357 19904
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12345 19867 12403 19873
rect 12710 19864 12716 19916
rect 12768 19864 12774 19916
rect 15286 19904 15292 19916
rect 12820 19876 15292 19904
rect 11425 19839 11483 19845
rect 11425 19836 11437 19839
rect 11072 19808 11437 19836
rect 11425 19805 11437 19808
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12728 19836 12756 19864
rect 12820 19845 12848 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15672 19904 15700 19944
rect 15746 19932 15752 19984
rect 15804 19972 15810 19984
rect 15804 19944 16436 19972
rect 15804 19932 15810 19944
rect 16408 19904 16436 19944
rect 19058 19932 19064 19984
rect 19116 19932 19122 19984
rect 19150 19932 19156 19984
rect 19208 19972 19214 19984
rect 19334 19972 19340 19984
rect 19208 19944 19340 19972
rect 19208 19932 19214 19944
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 19536 19904 19564 20012
rect 22094 20000 22100 20012
rect 22152 20040 22158 20052
rect 22281 20043 22339 20049
rect 22152 20012 22232 20040
rect 22152 20000 22158 20012
rect 21818 19972 21824 19984
rect 21376 19944 21824 19972
rect 15672 19876 16344 19904
rect 16408 19876 19564 19904
rect 12575 19808 12756 19836
rect 12805 19839 12863 19845
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12805 19805 12817 19839
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 13998 19796 14004 19848
rect 14056 19796 14062 19848
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16316 19845 16344 19876
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 21376 19904 21404 19944
rect 21818 19932 21824 19944
rect 21876 19932 21882 19984
rect 20956 19876 21404 19904
rect 20956 19864 20962 19876
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19836 16359 19839
rect 16669 19839 16727 19845
rect 16347 19808 16620 19836
rect 16347 19805 16359 19808
rect 16301 19799 16359 19805
rect 8312 19768 8340 19796
rect 11149 19771 11207 19777
rect 11149 19768 11161 19771
rect 8312 19740 11161 19768
rect 11149 19737 11161 19740
rect 11195 19737 11207 19771
rect 12713 19771 12771 19777
rect 11149 19731 11207 19737
rect 11256 19740 12434 19768
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 11256 19700 11284 19740
rect 1728 19672 11284 19700
rect 11609 19703 11667 19709
rect 1728 19660 1734 19672
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 11974 19700 11980 19712
rect 11655 19672 11980 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 12406 19700 12434 19740
rect 12713 19737 12725 19771
rect 12759 19768 12771 19771
rect 14016 19768 14044 19796
rect 12759 19740 14044 19768
rect 12759 19737 12771 19740
rect 12713 19731 12771 19737
rect 16022 19700 16028 19712
rect 12406 19672 16028 19700
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 16592 19700 16620 19808
rect 16669 19805 16681 19839
rect 16715 19836 16727 19839
rect 16758 19836 16764 19848
rect 16715 19808 16764 19836
rect 16715 19805 16727 19808
rect 16669 19799 16727 19805
rect 16758 19796 16764 19808
rect 16816 19836 16822 19848
rect 17402 19836 17408 19848
rect 16816 19808 17408 19836
rect 16816 19796 16822 19808
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 19334 19836 19340 19848
rect 18656 19808 19340 19836
rect 18656 19796 18662 19808
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19426 19796 19432 19848
rect 19484 19796 19490 19848
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19836 19763 19839
rect 19886 19836 19892 19848
rect 19751 19808 19892 19836
rect 19751 19805 19763 19808
rect 19705 19799 19763 19805
rect 19886 19796 19892 19808
rect 19944 19836 19950 19848
rect 19944 19808 20760 19836
rect 19944 19796 19950 19808
rect 20732 19780 20760 19808
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 20990 19836 20996 19848
rect 20864 19808 20996 19836
rect 20864 19796 20870 19808
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 21376 19845 21404 19876
rect 21450 19864 21456 19916
rect 21508 19904 21514 19916
rect 21612 19907 21670 19913
rect 21612 19904 21624 19907
rect 21508 19876 21624 19904
rect 21508 19864 21514 19876
rect 21612 19873 21624 19876
rect 21658 19904 21670 19907
rect 21658 19873 21680 19904
rect 21612 19867 21680 19873
rect 21361 19839 21419 19845
rect 21361 19805 21373 19839
rect 21407 19805 21419 19839
rect 21361 19799 21419 19805
rect 21652 19780 21680 19867
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 22097 19839 22155 19845
rect 22097 19836 22109 19839
rect 21784 19808 22109 19836
rect 21784 19796 21790 19808
rect 22097 19805 22109 19808
rect 22143 19805 22155 19839
rect 22204 19836 22232 20012
rect 22281 20009 22293 20043
rect 22327 20040 22339 20043
rect 22646 20040 22652 20052
rect 22327 20012 22652 20040
rect 22327 20009 22339 20012
rect 22281 20003 22339 20009
rect 22646 20000 22652 20012
rect 22704 20000 22710 20052
rect 22922 19972 22928 19984
rect 22756 19944 22928 19972
rect 22756 19904 22784 19944
rect 22922 19932 22928 19944
rect 22980 19972 22986 19984
rect 24394 19972 24400 19984
rect 22980 19944 24400 19972
rect 22980 19932 22986 19944
rect 24394 19932 24400 19944
rect 24452 19932 24458 19984
rect 24486 19932 24492 19984
rect 24544 19972 24550 19984
rect 24544 19944 26740 19972
rect 24544 19932 24550 19944
rect 22480 19876 22784 19904
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 22204 19808 22385 19836
rect 22097 19799 22155 19805
rect 22373 19805 22385 19808
rect 22419 19805 22431 19839
rect 22373 19799 22431 19805
rect 17494 19728 17500 19780
rect 17552 19768 17558 19780
rect 18693 19771 18751 19777
rect 18693 19768 18705 19771
rect 17552 19740 18705 19768
rect 17552 19728 17558 19740
rect 18693 19737 18705 19740
rect 18739 19737 18751 19771
rect 20254 19768 20260 19780
rect 18693 19731 18751 19737
rect 18800 19740 20260 19768
rect 18800 19700 18828 19740
rect 20254 19728 20260 19740
rect 20312 19728 20318 19780
rect 20349 19771 20407 19777
rect 20349 19737 20361 19771
rect 20395 19737 20407 19771
rect 20349 19731 20407 19737
rect 16592 19672 18828 19700
rect 18874 19660 18880 19712
rect 18932 19709 18938 19712
rect 18932 19703 18961 19709
rect 18949 19669 18961 19703
rect 18932 19663 18961 19669
rect 18932 19660 18938 19663
rect 19242 19660 19248 19712
rect 19300 19700 19306 19712
rect 19613 19703 19671 19709
rect 19613 19700 19625 19703
rect 19300 19672 19625 19700
rect 19300 19660 19306 19672
rect 19613 19669 19625 19672
rect 19659 19669 19671 19703
rect 20364 19700 20392 19731
rect 20438 19728 20444 19780
rect 20496 19728 20502 19780
rect 20714 19728 20720 19780
rect 20772 19728 20778 19780
rect 20901 19771 20959 19777
rect 20901 19737 20913 19771
rect 20947 19768 20959 19771
rect 21266 19768 21272 19780
rect 20947 19740 21272 19768
rect 20947 19737 20959 19740
rect 20901 19731 20959 19737
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 21542 19728 21548 19780
rect 21600 19728 21606 19780
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 22480 19768 22508 19876
rect 22646 19796 22652 19848
rect 22704 19796 22710 19848
rect 22756 19845 22784 19876
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19873 23443 19907
rect 23385 19867 23443 19873
rect 23860 19876 24624 19904
rect 22741 19839 22799 19845
rect 22741 19805 22753 19839
rect 22787 19805 22799 19839
rect 22741 19799 22799 19805
rect 23106 19796 23112 19848
rect 23164 19796 23170 19848
rect 21692 19740 22508 19768
rect 22664 19768 22692 19796
rect 23124 19768 23152 19796
rect 23400 19780 23428 19867
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 23658 19836 23664 19848
rect 23615 19808 23664 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 23658 19796 23664 19808
rect 23716 19796 23722 19848
rect 23860 19845 23888 19876
rect 23845 19839 23903 19845
rect 23845 19805 23857 19839
rect 23891 19805 23903 19839
rect 23845 19799 23903 19805
rect 23937 19839 23995 19845
rect 23937 19805 23949 19839
rect 23983 19805 23995 19839
rect 23937 19799 23995 19805
rect 22664 19740 23152 19768
rect 21692 19728 21698 19740
rect 23382 19728 23388 19780
rect 23440 19728 23446 19780
rect 23952 19768 23980 19799
rect 24026 19796 24032 19848
rect 24084 19836 24090 19848
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24084 19808 24409 19836
rect 24084 19796 24090 19808
rect 24397 19805 24409 19808
rect 24443 19836 24455 19839
rect 24486 19836 24492 19848
rect 24443 19808 24492 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 23492 19740 23980 19768
rect 21082 19700 21088 19712
rect 20364 19672 21088 19700
rect 19613 19663 19671 19669
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 21450 19660 21456 19712
rect 21508 19660 21514 19712
rect 21560 19700 21588 19728
rect 23492 19712 23520 19740
rect 21729 19703 21787 19709
rect 21729 19700 21741 19703
rect 21560 19672 21741 19700
rect 21729 19669 21741 19672
rect 21775 19669 21787 19703
rect 21729 19663 21787 19669
rect 21818 19660 21824 19712
rect 21876 19660 21882 19712
rect 21910 19660 21916 19712
rect 21968 19700 21974 19712
rect 22925 19703 22983 19709
rect 22925 19700 22937 19703
rect 21968 19672 22937 19700
rect 21968 19660 21974 19672
rect 22925 19669 22937 19672
rect 22971 19700 22983 19703
rect 23474 19700 23480 19712
rect 22971 19672 23480 19700
rect 22971 19669 22983 19672
rect 22925 19663 22983 19669
rect 23474 19660 23480 19672
rect 23532 19660 23538 19712
rect 24596 19709 24624 19876
rect 26712 19848 26740 19944
rect 26694 19796 26700 19848
rect 26752 19796 26758 19848
rect 24581 19703 24639 19709
rect 24581 19669 24593 19703
rect 24627 19700 24639 19703
rect 24762 19700 24768 19712
rect 24627 19672 24768 19700
rect 24627 19669 24639 19672
rect 24581 19663 24639 19669
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 26602 19660 26608 19712
rect 26660 19660 26666 19712
rect 1104 19610 31280 19632
rect 1104 19558 4922 19610
rect 4974 19558 4986 19610
rect 5038 19558 5050 19610
rect 5102 19558 5114 19610
rect 5166 19558 5178 19610
rect 5230 19558 5242 19610
rect 5294 19558 10922 19610
rect 10974 19558 10986 19610
rect 11038 19558 11050 19610
rect 11102 19558 11114 19610
rect 11166 19558 11178 19610
rect 11230 19558 11242 19610
rect 11294 19558 16922 19610
rect 16974 19558 16986 19610
rect 17038 19558 17050 19610
rect 17102 19558 17114 19610
rect 17166 19558 17178 19610
rect 17230 19558 17242 19610
rect 17294 19558 22922 19610
rect 22974 19558 22986 19610
rect 23038 19558 23050 19610
rect 23102 19558 23114 19610
rect 23166 19558 23178 19610
rect 23230 19558 23242 19610
rect 23294 19558 28922 19610
rect 28974 19558 28986 19610
rect 29038 19558 29050 19610
rect 29102 19558 29114 19610
rect 29166 19558 29178 19610
rect 29230 19558 29242 19610
rect 29294 19558 31280 19610
rect 1104 19536 31280 19558
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 14182 19496 14188 19508
rect 7616 19468 14188 19496
rect 7616 19456 7622 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 15286 19456 15292 19508
rect 15344 19496 15350 19508
rect 16117 19499 16175 19505
rect 16117 19496 16129 19499
rect 15344 19468 16129 19496
rect 15344 19456 15350 19468
rect 16117 19465 16129 19468
rect 16163 19465 16175 19499
rect 16117 19459 16175 19465
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 16482 19496 16488 19508
rect 16255 19468 16488 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 14826 19388 14832 19440
rect 14884 19428 14890 19440
rect 15473 19431 15531 19437
rect 15473 19428 15485 19431
rect 14884 19400 15485 19428
rect 14884 19388 14890 19400
rect 15473 19397 15485 19400
rect 15519 19428 15531 19431
rect 15746 19428 15752 19440
rect 15519 19400 15752 19428
rect 15519 19397 15531 19400
rect 15473 19391 15531 19397
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 15838 19388 15844 19440
rect 15896 19388 15902 19440
rect 16132 19428 16160 19459
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 22554 19496 22560 19508
rect 19208 19468 22560 19496
rect 19208 19456 19214 19468
rect 22554 19456 22560 19468
rect 22612 19496 22618 19508
rect 23750 19496 23756 19508
rect 22612 19468 23756 19496
rect 22612 19456 22618 19468
rect 23750 19456 23756 19468
rect 23808 19456 23814 19508
rect 26789 19499 26847 19505
rect 26789 19496 26801 19499
rect 24964 19468 26801 19496
rect 19168 19428 19196 19456
rect 16132 19400 19196 19428
rect 19242 19388 19248 19440
rect 19300 19428 19306 19440
rect 20073 19431 20131 19437
rect 19300 19388 19334 19428
rect 20073 19397 20085 19431
rect 20119 19428 20131 19431
rect 21450 19428 21456 19440
rect 20119 19400 21456 19428
rect 20119 19397 20131 19400
rect 20073 19391 20131 19397
rect 21450 19388 21456 19400
rect 21508 19388 21514 19440
rect 2777 19363 2835 19369
rect 2777 19329 2789 19363
rect 2823 19360 2835 19363
rect 3326 19360 3332 19372
rect 2823 19332 3332 19360
rect 2823 19329 2835 19332
rect 2777 19323 2835 19329
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 15289 19363 15347 19369
rect 15289 19329 15301 19363
rect 15335 19360 15347 19363
rect 15562 19360 15568 19372
rect 15335 19332 15568 19360
rect 15335 19329 15347 19332
rect 15289 19323 15347 19329
rect 15562 19320 15568 19332
rect 15620 19320 15626 19372
rect 15856 19360 15884 19388
rect 17313 19363 17371 19369
rect 17313 19360 17325 19363
rect 15856 19332 17325 19360
rect 17313 19329 17325 19332
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 17402 19320 17408 19372
rect 17460 19320 17466 19372
rect 17678 19320 17684 19372
rect 17736 19320 17742 19372
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19329 17923 19363
rect 19306 19360 19334 19388
rect 24964 19372 24992 19468
rect 26789 19465 26801 19468
rect 26835 19465 26847 19499
rect 26789 19459 26847 19465
rect 26602 19428 26608 19440
rect 26542 19400 26608 19428
rect 26602 19388 26608 19400
rect 26660 19388 26666 19440
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19306 19332 19441 19360
rect 17865 19323 17923 19329
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4614 19292 4620 19304
rect 4479 19264 4620 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 5074 19252 5080 19304
rect 5132 19292 5138 19304
rect 16393 19295 16451 19301
rect 5132 19264 15884 19292
rect 5132 19252 5138 19264
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 15749 19227 15807 19233
rect 15749 19224 15761 19227
rect 15252 19196 15761 19224
rect 15252 19184 15258 19196
rect 15749 19193 15761 19196
rect 15795 19193 15807 19227
rect 15856 19224 15884 19264
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 16574 19292 16580 19304
rect 16439 19264 16580 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19292 17003 19295
rect 17221 19295 17279 19301
rect 16991 19264 17080 19292
rect 16991 19261 17003 19264
rect 16945 19255 17003 19261
rect 17052 19224 17080 19264
rect 17221 19261 17233 19295
rect 17267 19292 17279 19295
rect 17420 19292 17448 19320
rect 17267 19264 17448 19292
rect 17880 19292 17908 19323
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 20438 19360 20444 19372
rect 19904 19332 20444 19360
rect 19797 19295 19855 19301
rect 19797 19292 19809 19295
rect 17880 19264 19809 19292
rect 17267 19261 17279 19264
rect 17221 19255 17279 19261
rect 15856 19196 17080 19224
rect 15749 19187 15807 19193
rect 2590 19116 2596 19168
rect 2648 19116 2654 19168
rect 3786 19116 3792 19168
rect 3844 19116 3850 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4706 19156 4712 19168
rect 4120 19128 4712 19156
rect 4120 19116 4126 19128
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 15470 19156 15476 19168
rect 10100 19128 15476 19156
rect 10100 19116 10106 19128
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15654 19116 15660 19168
rect 15712 19116 15718 19168
rect 17052 19156 17080 19196
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 17880 19224 17908 19264
rect 19797 19261 19809 19264
rect 19843 19261 19855 19295
rect 19797 19255 19855 19261
rect 17368 19196 17908 19224
rect 17368 19184 17374 19196
rect 18230 19184 18236 19236
rect 18288 19224 18294 19236
rect 18598 19224 18604 19236
rect 18288 19196 18604 19224
rect 18288 19184 18294 19196
rect 18598 19184 18604 19196
rect 18656 19224 18662 19236
rect 19904 19224 19932 19332
rect 20438 19320 20444 19332
rect 20496 19320 20502 19372
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20898 19360 20904 19372
rect 20579 19332 20904 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 20990 19320 20996 19372
rect 21048 19320 21054 19372
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 22094 19360 22100 19372
rect 21140 19332 22100 19360
rect 21140 19320 21146 19332
rect 22094 19320 22100 19332
rect 22152 19360 22158 19372
rect 22646 19360 22652 19372
rect 22152 19332 22652 19360
rect 22152 19320 22158 19332
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 24946 19320 24952 19372
rect 25004 19320 25010 19372
rect 25038 19320 25044 19372
rect 25096 19320 25102 19372
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 30561 19363 30619 19369
rect 30561 19360 30573 19363
rect 29696 19332 30573 19360
rect 29696 19320 29702 19332
rect 30561 19329 30573 19332
rect 30607 19329 30619 19363
rect 30561 19323 30619 19329
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 21174 19292 21180 19304
rect 20680 19264 21180 19292
rect 20680 19252 20686 19264
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21266 19252 21272 19304
rect 21324 19292 21330 19304
rect 21545 19295 21603 19301
rect 21545 19292 21557 19295
rect 21324 19264 21557 19292
rect 21324 19252 21330 19264
rect 21545 19261 21557 19264
rect 21591 19292 21603 19295
rect 21910 19292 21916 19304
rect 21591 19264 21916 19292
rect 21591 19261 21603 19264
rect 21545 19255 21603 19261
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 18656 19196 19932 19224
rect 18656 19184 18662 19196
rect 17586 19156 17592 19168
rect 17052 19128 17592 19156
rect 17586 19116 17592 19128
rect 17644 19116 17650 19168
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19521 19159 19579 19165
rect 19521 19156 19533 19159
rect 18932 19128 19533 19156
rect 18932 19116 18938 19128
rect 19521 19125 19533 19128
rect 19567 19125 19579 19159
rect 19521 19119 19579 19125
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 23474 19156 23480 19168
rect 21600 19128 23480 19156
rect 21600 19116 21606 19128
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 24394 19116 24400 19168
rect 24452 19156 24458 19168
rect 24765 19159 24823 19165
rect 24765 19156 24777 19159
rect 24452 19128 24777 19156
rect 24452 19116 24458 19128
rect 24765 19125 24777 19128
rect 24811 19125 24823 19159
rect 24765 19119 24823 19125
rect 30837 19159 30895 19165
rect 30837 19125 30849 19159
rect 30883 19156 30895 19159
rect 30926 19156 30932 19168
rect 30883 19128 30932 19156
rect 30883 19125 30895 19128
rect 30837 19119 30895 19125
rect 30926 19116 30932 19128
rect 30984 19116 30990 19168
rect 1104 19066 31280 19088
rect 1104 19014 4182 19066
rect 4234 19014 4246 19066
rect 4298 19014 4310 19066
rect 4362 19014 4374 19066
rect 4426 19014 4438 19066
rect 4490 19014 4502 19066
rect 4554 19014 10182 19066
rect 10234 19014 10246 19066
rect 10298 19014 10310 19066
rect 10362 19014 10374 19066
rect 10426 19014 10438 19066
rect 10490 19014 10502 19066
rect 10554 19014 16182 19066
rect 16234 19014 16246 19066
rect 16298 19014 16310 19066
rect 16362 19014 16374 19066
rect 16426 19014 16438 19066
rect 16490 19014 16502 19066
rect 16554 19014 22182 19066
rect 22234 19014 22246 19066
rect 22298 19014 22310 19066
rect 22362 19014 22374 19066
rect 22426 19014 22438 19066
rect 22490 19014 22502 19066
rect 22554 19014 28182 19066
rect 28234 19014 28246 19066
rect 28298 19014 28310 19066
rect 28362 19014 28374 19066
rect 28426 19014 28438 19066
rect 28490 19014 28502 19066
rect 28554 19014 31280 19066
rect 1104 18992 31280 19014
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3384 18924 3801 18952
rect 3384 18912 3390 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 4580 18924 5304 18952
rect 4580 18912 4586 18924
rect 3605 18887 3663 18893
rect 3605 18853 3617 18887
rect 3651 18884 3663 18887
rect 4706 18884 4712 18896
rect 3651 18856 4712 18884
rect 3651 18853 3663 18856
rect 3605 18847 3663 18853
rect 4706 18844 4712 18856
rect 4764 18884 4770 18896
rect 5276 18884 5304 18924
rect 6546 18912 6552 18964
rect 6604 18952 6610 18964
rect 6917 18955 6975 18961
rect 6917 18952 6929 18955
rect 6604 18924 6929 18952
rect 6604 18912 6610 18924
rect 6917 18921 6929 18924
rect 6963 18921 6975 18955
rect 16298 18952 16304 18964
rect 6917 18915 6975 18921
rect 9646 18924 16304 18952
rect 9646 18884 9674 18924
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 19794 18952 19800 18964
rect 16408 18924 19800 18952
rect 4764 18856 5212 18884
rect 5276 18856 9674 18884
rect 14553 18887 14611 18893
rect 4764 18844 4770 18856
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 4028 18788 4445 18816
rect 4028 18776 4034 18788
rect 4433 18785 4445 18788
rect 4479 18816 4491 18819
rect 5074 18816 5080 18828
rect 4479 18788 5080 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 5074 18776 5080 18788
rect 5132 18776 5138 18828
rect 5184 18825 5212 18856
rect 14553 18853 14565 18887
rect 14599 18884 14611 18887
rect 15102 18884 15108 18896
rect 14599 18856 15108 18884
rect 14599 18853 14611 18856
rect 14553 18847 14611 18853
rect 15102 18844 15108 18856
rect 15160 18844 15166 18896
rect 16408 18884 16436 18924
rect 19794 18912 19800 18924
rect 19852 18912 19858 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 20916 18924 21465 18952
rect 15580 18856 16436 18884
rect 16500 18856 17448 18884
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18785 5227 18819
rect 15580 18816 15608 18856
rect 16500 18828 16528 18856
rect 17420 18828 17448 18856
rect 5169 18779 5227 18785
rect 6748 18788 9812 18816
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 4798 18748 4804 18760
rect 2280 18720 4804 18748
rect 2280 18708 2286 18720
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 6748 18757 6776 18788
rect 9784 18760 9812 18788
rect 12406 18788 15608 18816
rect 6733 18751 6791 18757
rect 6733 18717 6745 18751
rect 6779 18717 6791 18751
rect 6733 18711 6791 18717
rect 2492 18683 2550 18689
rect 2492 18649 2504 18683
rect 2538 18680 2550 18683
rect 2590 18680 2596 18692
rect 2538 18652 2596 18680
rect 2538 18649 2550 18652
rect 2492 18643 2550 18649
rect 2590 18640 2596 18652
rect 2648 18640 2654 18692
rect 4157 18683 4215 18689
rect 4157 18649 4169 18683
rect 4203 18680 4215 18683
rect 4617 18683 4675 18689
rect 4617 18680 4629 18683
rect 4203 18652 4629 18680
rect 4203 18649 4215 18652
rect 4157 18643 4215 18649
rect 4617 18649 4629 18652
rect 4663 18649 4675 18683
rect 4617 18643 4675 18649
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 6454 18612 6460 18624
rect 4304 18584 6460 18612
rect 4304 18572 4310 18584
rect 6454 18572 6460 18584
rect 6512 18612 6518 18624
rect 6748 18612 6776 18711
rect 9306 18708 9312 18760
rect 9364 18708 9370 18760
rect 9766 18708 9772 18760
rect 9824 18708 9830 18760
rect 6822 18640 6828 18692
rect 6880 18680 6886 18692
rect 12406 18680 12434 18788
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18748 12955 18751
rect 14090 18748 14096 18760
rect 12943 18720 14096 18748
rect 12943 18717 12955 18720
rect 12897 18711 12955 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 14734 18748 14740 18760
rect 14240 18720 14740 18748
rect 14240 18708 14246 18720
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 6880 18652 12434 18680
rect 15580 18680 15608 18788
rect 15654 18776 15660 18828
rect 15712 18776 15718 18828
rect 16482 18776 16488 18828
rect 16540 18776 16546 18828
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 17402 18776 17408 18828
rect 17460 18776 17466 18828
rect 17494 18776 17500 18828
rect 17552 18816 17558 18828
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 17552 18788 17601 18816
rect 17552 18776 17558 18788
rect 17589 18785 17601 18788
rect 17635 18785 17647 18819
rect 17589 18779 17647 18785
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 20717 18819 20775 18825
rect 20717 18816 20729 18819
rect 18012 18788 20729 18816
rect 18012 18776 18018 18788
rect 20717 18785 20729 18788
rect 20763 18785 20775 18819
rect 20717 18779 20775 18785
rect 15672 18748 15700 18776
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15672 18720 16405 18748
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 17681 18751 17739 18757
rect 16816 18720 17540 18748
rect 16816 18708 16822 18720
rect 15749 18683 15807 18689
rect 15749 18680 15761 18683
rect 15580 18652 15761 18680
rect 6880 18640 6886 18652
rect 15749 18649 15761 18652
rect 15795 18649 15807 18683
rect 15749 18643 15807 18649
rect 17037 18683 17095 18689
rect 17037 18649 17049 18683
rect 17083 18680 17095 18683
rect 17402 18680 17408 18692
rect 17083 18652 17408 18680
rect 17083 18649 17095 18652
rect 17037 18643 17095 18649
rect 17402 18640 17408 18652
rect 17460 18640 17466 18692
rect 17512 18680 17540 18720
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 17862 18748 17868 18760
rect 17727 18720 17868 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 19702 18748 19708 18760
rect 18279 18720 19708 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18064 18680 18092 18711
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 17512 18652 18092 18680
rect 20916 18680 20944 18924
rect 21453 18921 21465 18924
rect 21499 18952 21511 18955
rect 21726 18952 21732 18964
rect 21499 18924 21732 18952
rect 21499 18921 21511 18924
rect 21453 18915 21511 18921
rect 21726 18912 21732 18924
rect 21784 18912 21790 18964
rect 24486 18912 24492 18964
rect 24544 18912 24550 18964
rect 25314 18912 25320 18964
rect 25372 18912 25378 18964
rect 21818 18884 21824 18896
rect 21008 18856 21824 18884
rect 21008 18757 21036 18856
rect 21818 18844 21824 18856
rect 21876 18884 21882 18896
rect 23566 18884 23572 18896
rect 21876 18856 23572 18884
rect 21876 18844 21882 18856
rect 21634 18776 21640 18828
rect 21692 18776 21698 18828
rect 22020 18825 22048 18856
rect 23566 18844 23572 18856
rect 23624 18884 23630 18896
rect 24670 18884 24676 18896
rect 23624 18856 24676 18884
rect 23624 18844 23630 18856
rect 24670 18844 24676 18856
rect 24728 18884 24734 18896
rect 24765 18887 24823 18893
rect 24765 18884 24777 18887
rect 24728 18856 24777 18884
rect 24728 18844 24734 18856
rect 24765 18853 24777 18856
rect 24811 18853 24823 18887
rect 24765 18847 24823 18853
rect 22005 18819 22063 18825
rect 22005 18785 22017 18819
rect 22051 18816 22063 18819
rect 22051 18788 22085 18816
rect 22051 18785 22063 18788
rect 22005 18779 22063 18785
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18717 21051 18751
rect 20993 18711 21051 18717
rect 21542 18708 21548 18760
rect 21600 18708 21606 18760
rect 25130 18708 25136 18760
rect 25188 18708 25194 18760
rect 21085 18683 21143 18689
rect 21085 18680 21097 18683
rect 20916 18652 21097 18680
rect 17696 18624 17724 18652
rect 21085 18649 21097 18652
rect 21131 18649 21143 18683
rect 21085 18643 21143 18649
rect 21266 18640 21272 18692
rect 21324 18640 21330 18692
rect 6512 18584 6776 18612
rect 6512 18572 6518 18584
rect 9122 18572 9128 18624
rect 9180 18572 9186 18624
rect 12710 18572 12716 18624
rect 12768 18572 12774 18624
rect 17678 18572 17684 18624
rect 17736 18572 17742 18624
rect 20901 18615 20959 18621
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21560 18612 21588 18708
rect 24581 18683 24639 18689
rect 24581 18649 24593 18683
rect 24627 18680 24639 18683
rect 24949 18683 25007 18689
rect 24949 18680 24961 18683
rect 24627 18652 24716 18680
rect 24627 18649 24639 18652
rect 24581 18643 24639 18649
rect 24688 18624 24716 18652
rect 24872 18652 24961 18680
rect 24872 18624 24900 18652
rect 24949 18649 24961 18652
rect 24995 18649 25007 18683
rect 24949 18643 25007 18649
rect 20947 18584 21588 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21818 18572 21824 18624
rect 21876 18572 21882 18624
rect 24670 18572 24676 18624
rect 24728 18572 24734 18624
rect 24854 18572 24860 18624
rect 24912 18572 24918 18624
rect 1104 18522 31280 18544
rect 1104 18470 4922 18522
rect 4974 18470 4986 18522
rect 5038 18470 5050 18522
rect 5102 18470 5114 18522
rect 5166 18470 5178 18522
rect 5230 18470 5242 18522
rect 5294 18470 10922 18522
rect 10974 18470 10986 18522
rect 11038 18470 11050 18522
rect 11102 18470 11114 18522
rect 11166 18470 11178 18522
rect 11230 18470 11242 18522
rect 11294 18470 16922 18522
rect 16974 18470 16986 18522
rect 17038 18470 17050 18522
rect 17102 18470 17114 18522
rect 17166 18470 17178 18522
rect 17230 18470 17242 18522
rect 17294 18470 22922 18522
rect 22974 18470 22986 18522
rect 23038 18470 23050 18522
rect 23102 18470 23114 18522
rect 23166 18470 23178 18522
rect 23230 18470 23242 18522
rect 23294 18470 28922 18522
rect 28974 18470 28986 18522
rect 29038 18470 29050 18522
rect 29102 18470 29114 18522
rect 29166 18470 29178 18522
rect 29230 18470 29242 18522
rect 29294 18470 31280 18522
rect 1104 18448 31280 18470
rect 2222 18368 2228 18420
rect 2280 18368 2286 18420
rect 3513 18411 3571 18417
rect 3513 18377 3525 18411
rect 3559 18377 3571 18411
rect 3513 18371 3571 18377
rect 1394 18232 1400 18284
rect 1452 18232 1458 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2240 18272 2268 18368
rect 3528 18340 3556 18371
rect 3786 18368 3792 18420
rect 3844 18408 3850 18420
rect 3973 18411 4031 18417
rect 3973 18408 3985 18411
rect 3844 18380 3985 18408
rect 3844 18368 3850 18380
rect 3973 18377 3985 18380
rect 4019 18377 4031 18411
rect 3973 18371 4031 18377
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18408 4123 18411
rect 4246 18408 4252 18420
rect 4111 18380 4252 18408
rect 4111 18377 4123 18380
rect 4065 18371 4123 18377
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 4614 18408 4620 18420
rect 4448 18380 4620 18408
rect 4448 18340 4476 18380
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 4706 18368 4712 18420
rect 4764 18368 4770 18420
rect 6365 18411 6423 18417
rect 6365 18377 6377 18411
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 3528 18312 4476 18340
rect 2406 18281 2412 18284
rect 2179 18244 2268 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2400 18235 2412 18281
rect 2406 18232 2412 18235
rect 2464 18232 2470 18284
rect 4448 18281 4476 18312
rect 4522 18300 4528 18352
rect 4580 18300 4586 18352
rect 4433 18275 4491 18281
rect 4433 18241 4445 18275
rect 4479 18241 4491 18275
rect 4540 18272 4568 18300
rect 4724 18281 4752 18368
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 4540 18244 4629 18272
rect 4433 18235 4491 18241
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 5442 18272 5448 18284
rect 4847 18244 5448 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 6089 18275 6147 18281
rect 6089 18241 6101 18275
rect 6135 18272 6147 18275
rect 6380 18272 6408 18371
rect 6546 18368 6552 18420
rect 6604 18408 6610 18420
rect 6730 18408 6736 18420
rect 6604 18380 6736 18408
rect 6604 18368 6610 18380
rect 6730 18368 6736 18380
rect 6788 18408 6794 18420
rect 6825 18411 6883 18417
rect 6825 18408 6837 18411
rect 6788 18380 6837 18408
rect 6788 18368 6794 18380
rect 6825 18377 6837 18380
rect 6871 18408 6883 18411
rect 6871 18380 8984 18408
rect 6871 18377 6883 18380
rect 6825 18371 6883 18377
rect 6135 18244 6408 18272
rect 6472 18312 7328 18340
rect 6135 18241 6147 18244
rect 6089 18235 6147 18241
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 3292 18176 4261 18204
rect 3292 18164 3298 18176
rect 4249 18173 4261 18176
rect 4295 18204 4307 18207
rect 6472 18204 6500 18312
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 6779 18244 7205 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 4295 18176 6500 18204
rect 4295 18173 4307 18176
rect 4249 18167 4307 18173
rect 6822 18164 6828 18216
rect 6880 18204 6886 18216
rect 6917 18207 6975 18213
rect 6917 18204 6929 18207
rect 6880 18176 6929 18204
rect 6880 18164 6886 18176
rect 6917 18173 6929 18176
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 4985 18139 5043 18145
rect 3528 18108 4108 18136
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 3050 18068 3056 18080
rect 1627 18040 3056 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 3050 18028 3056 18040
rect 3108 18068 3114 18080
rect 3528 18068 3556 18108
rect 4080 18080 4108 18108
rect 4985 18105 4997 18139
rect 5031 18136 5043 18139
rect 6454 18136 6460 18148
rect 5031 18108 6460 18136
rect 5031 18105 5043 18108
rect 4985 18099 5043 18105
rect 6454 18096 6460 18108
rect 6512 18096 6518 18148
rect 3108 18040 3556 18068
rect 3108 18028 3114 18040
rect 3602 18028 3608 18080
rect 3660 18028 3666 18080
rect 4062 18028 4068 18080
rect 4120 18028 4126 18080
rect 5902 18028 5908 18080
rect 5960 18028 5966 18080
rect 7300 18068 7328 18312
rect 8386 18300 8392 18352
rect 8444 18300 8450 18352
rect 8018 18232 8024 18284
rect 8076 18232 8082 18284
rect 8956 18272 8984 18380
rect 9122 18368 9128 18420
rect 9180 18368 9186 18420
rect 10137 18411 10195 18417
rect 10137 18377 10149 18411
rect 10183 18377 10195 18411
rect 10137 18371 10195 18377
rect 15749 18411 15807 18417
rect 15749 18377 15761 18411
rect 15795 18408 15807 18411
rect 15930 18408 15936 18420
rect 15795 18380 15936 18408
rect 15795 18377 15807 18380
rect 15749 18371 15807 18377
rect 9024 18343 9082 18349
rect 9024 18309 9036 18343
rect 9070 18340 9082 18343
rect 9140 18340 9168 18368
rect 9070 18312 9168 18340
rect 9070 18309 9082 18312
rect 9024 18303 9082 18309
rect 10152 18272 10180 18371
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 16724 18380 18061 18408
rect 16724 18368 16730 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 23753 18411 23811 18417
rect 23753 18408 23765 18411
rect 18049 18371 18107 18377
rect 23492 18380 23765 18408
rect 23492 18352 23520 18380
rect 23753 18377 23765 18380
rect 23799 18377 23811 18411
rect 25317 18411 25375 18417
rect 25317 18408 25329 18411
rect 23753 18371 23811 18377
rect 23860 18380 25329 18408
rect 12710 18349 12716 18352
rect 12693 18343 12716 18349
rect 12693 18309 12705 18343
rect 12693 18303 12716 18309
rect 12710 18300 12716 18303
rect 12768 18300 12774 18352
rect 15838 18300 15844 18352
rect 15896 18340 15902 18352
rect 16117 18343 16175 18349
rect 16117 18340 16129 18343
rect 15896 18312 16129 18340
rect 15896 18300 15902 18312
rect 16117 18309 16129 18312
rect 16163 18309 16175 18343
rect 16482 18340 16488 18352
rect 16117 18303 16175 18309
rect 16224 18312 16488 18340
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 8956 18244 10088 18272
rect 10152 18244 10793 18272
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 8110 18204 8116 18216
rect 7883 18176 8116 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 10060 18204 10088 18244
rect 10781 18241 10793 18244
rect 10827 18272 10839 18275
rect 11606 18272 11612 18284
rect 10827 18244 11612 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 11606 18232 11612 18244
rect 11664 18232 11670 18284
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18272 15163 18275
rect 15194 18272 15200 18284
rect 15151 18244 15200 18272
rect 15151 18241 15163 18244
rect 15105 18235 15163 18241
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16022 18272 16028 18284
rect 15703 18244 16028 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16022 18232 16028 18244
rect 16080 18272 16086 18284
rect 16224 18272 16252 18312
rect 16482 18300 16488 18312
rect 16540 18340 16546 18352
rect 16758 18340 16764 18352
rect 16540 18312 16764 18340
rect 16540 18300 16546 18312
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 18141 18343 18199 18349
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 18414 18340 18420 18352
rect 18187 18312 18420 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 18414 18300 18420 18312
rect 18472 18340 18478 18352
rect 23382 18340 23388 18352
rect 18472 18312 23388 18340
rect 18472 18300 18478 18312
rect 23382 18300 23388 18312
rect 23440 18300 23446 18352
rect 23474 18300 23480 18352
rect 23532 18300 23538 18352
rect 23566 18300 23572 18352
rect 23624 18300 23630 18352
rect 16080 18244 16252 18272
rect 16080 18232 16086 18244
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16356 18244 16681 18272
rect 16356 18232 16362 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16850 18232 16856 18284
rect 16908 18232 16914 18284
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19242 18272 19248 18284
rect 19024 18244 19248 18272
rect 19024 18232 19030 18244
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19429 18275 19487 18281
rect 19429 18241 19441 18275
rect 19475 18272 19487 18275
rect 19702 18272 19708 18284
rect 19475 18244 19708 18272
rect 19475 18241 19487 18244
rect 19429 18235 19487 18241
rect 10594 18204 10600 18216
rect 10060 18176 10600 18204
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 14274 18164 14280 18216
rect 14332 18164 14338 18216
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18204 15347 18207
rect 15470 18204 15476 18216
rect 15335 18176 15476 18204
rect 15335 18173 15347 18176
rect 15289 18167 15347 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 15988 18176 16221 18204
rect 15988 18164 15994 18176
rect 16209 18173 16221 18176
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 16393 18207 16451 18213
rect 16393 18173 16405 18207
rect 16439 18204 16451 18207
rect 16574 18204 16580 18216
rect 16439 18176 16580 18204
rect 16439 18173 16451 18176
rect 16393 18167 16451 18173
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 17313 18207 17371 18213
rect 17313 18173 17325 18207
rect 17359 18204 17371 18207
rect 17494 18204 17500 18216
rect 17359 18176 17500 18204
rect 17359 18173 17371 18176
rect 17313 18167 17371 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 17589 18207 17647 18213
rect 17589 18173 17601 18207
rect 17635 18204 17647 18207
rect 17770 18204 17776 18216
rect 17635 18176 17776 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 9950 18096 9956 18148
rect 10008 18136 10014 18148
rect 10229 18139 10287 18145
rect 10229 18136 10241 18139
rect 10008 18108 10241 18136
rect 10008 18096 10014 18108
rect 10229 18105 10241 18108
rect 10275 18105 10287 18139
rect 10229 18099 10287 18105
rect 13817 18139 13875 18145
rect 13817 18105 13829 18139
rect 13863 18136 13875 18139
rect 14292 18136 14320 18164
rect 17604 18136 17632 18167
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 19444 18136 19472 18235
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18272 21327 18275
rect 21542 18272 21548 18284
rect 21315 18244 21548 18272
rect 21315 18241 21327 18244
rect 21269 18235 21327 18241
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23584 18272 23612 18300
rect 23339 18244 23612 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 23860 18204 23888 18380
rect 25317 18377 25329 18380
rect 25363 18377 25375 18411
rect 25317 18371 25375 18377
rect 24394 18300 24400 18352
rect 24452 18300 24458 18352
rect 23934 18232 23940 18284
rect 23992 18272 23998 18284
rect 24029 18275 24087 18281
rect 24029 18272 24041 18275
rect 23992 18244 24041 18272
rect 23992 18232 23998 18244
rect 24029 18241 24041 18244
rect 24075 18272 24087 18275
rect 24673 18275 24731 18281
rect 24673 18272 24685 18275
rect 24075 18244 24685 18272
rect 24075 18241 24087 18244
rect 24029 18235 24087 18241
rect 24673 18241 24685 18244
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 24946 18232 24952 18284
rect 25004 18232 25010 18284
rect 27065 18275 27123 18281
rect 27065 18241 27077 18275
rect 27111 18241 27123 18275
rect 27065 18235 27123 18241
rect 20772 18176 23888 18204
rect 24213 18207 24271 18213
rect 20772 18164 20778 18176
rect 24213 18173 24225 18207
rect 24259 18173 24271 18207
rect 24964 18204 24992 18232
rect 25041 18207 25099 18213
rect 25041 18204 25053 18207
rect 24964 18176 25053 18204
rect 24213 18167 24271 18173
rect 25041 18173 25053 18176
rect 25087 18173 25099 18207
rect 25041 18167 25099 18173
rect 13863 18108 14320 18136
rect 14476 18108 17632 18136
rect 17696 18108 19472 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 14476 18068 14504 18108
rect 7300 18040 14504 18068
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 14829 18071 14887 18077
rect 14829 18068 14841 18071
rect 14608 18040 14841 18068
rect 14608 18028 14614 18040
rect 14829 18037 14841 18040
rect 14875 18037 14887 18071
rect 14829 18031 14887 18037
rect 15102 18028 15108 18080
rect 15160 18068 15166 18080
rect 17696 18068 17724 18108
rect 19610 18096 19616 18148
rect 19668 18136 19674 18148
rect 24228 18136 24256 18167
rect 26694 18164 26700 18216
rect 26752 18204 26758 18216
rect 26970 18204 26976 18216
rect 26752 18176 26976 18204
rect 26752 18164 26758 18176
rect 26970 18164 26976 18176
rect 27028 18204 27034 18216
rect 27080 18204 27108 18235
rect 27028 18176 27108 18204
rect 27028 18164 27034 18176
rect 24854 18145 24860 18148
rect 24838 18139 24860 18145
rect 24838 18136 24850 18139
rect 19668 18108 21312 18136
rect 24228 18108 24850 18136
rect 19668 18096 19674 18108
rect 21284 18080 21312 18108
rect 24838 18105 24850 18108
rect 24912 18136 24918 18148
rect 24912 18108 27660 18136
rect 24838 18099 24860 18105
rect 24854 18096 24860 18099
rect 24912 18096 24918 18108
rect 27632 18080 27660 18108
rect 15160 18040 17724 18068
rect 19429 18071 19487 18077
rect 15160 18028 15166 18040
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 20070 18068 20076 18080
rect 19475 18040 20076 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 21266 18028 21272 18080
rect 21324 18028 21330 18080
rect 21358 18028 21364 18080
rect 21416 18028 21422 18080
rect 23106 18028 23112 18080
rect 23164 18028 23170 18080
rect 24026 18028 24032 18080
rect 24084 18028 24090 18080
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 24670 18068 24676 18080
rect 24351 18040 24676 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 24670 18028 24676 18040
rect 24728 18068 24734 18080
rect 24949 18071 25007 18077
rect 24949 18068 24961 18071
rect 24728 18040 24961 18068
rect 24728 18028 24734 18040
rect 24949 18037 24961 18040
rect 24995 18068 25007 18071
rect 26326 18068 26332 18080
rect 24995 18040 26332 18068
rect 24995 18037 25007 18040
rect 24949 18031 25007 18037
rect 26326 18028 26332 18040
rect 26384 18028 26390 18080
rect 27062 18028 27068 18080
rect 27120 18068 27126 18080
rect 27157 18071 27215 18077
rect 27157 18068 27169 18071
rect 27120 18040 27169 18068
rect 27120 18028 27126 18040
rect 27157 18037 27169 18040
rect 27203 18037 27215 18071
rect 27157 18031 27215 18037
rect 27614 18028 27620 18080
rect 27672 18028 27678 18080
rect 1104 17978 31280 18000
rect 1104 17926 4182 17978
rect 4234 17926 4246 17978
rect 4298 17926 4310 17978
rect 4362 17926 4374 17978
rect 4426 17926 4438 17978
rect 4490 17926 4502 17978
rect 4554 17926 10182 17978
rect 10234 17926 10246 17978
rect 10298 17926 10310 17978
rect 10362 17926 10374 17978
rect 10426 17926 10438 17978
rect 10490 17926 10502 17978
rect 10554 17926 16182 17978
rect 16234 17926 16246 17978
rect 16298 17926 16310 17978
rect 16362 17926 16374 17978
rect 16426 17926 16438 17978
rect 16490 17926 16502 17978
rect 16554 17926 22182 17978
rect 22234 17926 22246 17978
rect 22298 17926 22310 17978
rect 22362 17926 22374 17978
rect 22426 17926 22438 17978
rect 22490 17926 22502 17978
rect 22554 17926 28182 17978
rect 28234 17926 28246 17978
rect 28298 17926 28310 17978
rect 28362 17926 28374 17978
rect 28426 17926 28438 17978
rect 28490 17926 28502 17978
rect 28554 17926 31280 17978
rect 1104 17904 31280 17926
rect 2406 17824 2412 17876
rect 2464 17864 2470 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 2464 17836 2513 17864
rect 2464 17824 2470 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 2501 17827 2559 17833
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 5500 17836 7972 17864
rect 5500 17824 5506 17836
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 4856 17700 5457 17728
rect 4856 17688 4862 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 7944 17728 7972 17836
rect 9306 17824 9312 17876
rect 9364 17824 9370 17876
rect 12250 17864 12256 17876
rect 9416 17836 12256 17864
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 9416 17796 9444 17836
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 12406 17836 13676 17864
rect 8260 17768 9444 17796
rect 8260 17756 8266 17768
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 12406 17796 12434 17836
rect 9732 17768 12434 17796
rect 9732 17756 9738 17768
rect 9582 17728 9588 17740
rect 7944 17700 9588 17728
rect 5445 17691 5503 17697
rect 2685 17663 2743 17669
rect 2685 17629 2697 17663
rect 2731 17660 2743 17663
rect 3602 17660 3608 17672
rect 2731 17632 3608 17660
rect 2731 17629 2743 17632
rect 2685 17623 2743 17629
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 5460 17660 5488 17691
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 9876 17737 9904 17768
rect 13648 17740 13676 17836
rect 14090 17824 14096 17876
rect 14148 17824 14154 17876
rect 16025 17867 16083 17873
rect 16025 17833 16037 17867
rect 16071 17864 16083 17867
rect 17218 17864 17224 17876
rect 16071 17836 17224 17864
rect 16071 17833 16083 17836
rect 16025 17827 16083 17833
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 18877 17867 18935 17873
rect 18877 17864 18889 17867
rect 18524 17836 18889 17864
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15930 17796 15936 17808
rect 15252 17768 15936 17796
rect 15252 17756 15258 17768
rect 15930 17756 15936 17768
rect 15988 17796 15994 17808
rect 16850 17796 16856 17808
rect 15988 17768 16160 17796
rect 15988 17756 15994 17768
rect 9861 17731 9919 17737
rect 9861 17697 9873 17731
rect 9907 17697 9919 17731
rect 11882 17728 11888 17740
rect 9861 17691 9919 17697
rect 11348 17700 11888 17728
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 5460 17632 6929 17660
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17660 9735 17663
rect 9950 17660 9956 17672
rect 9723 17632 9956 17660
rect 9723 17629 9735 17632
rect 9677 17623 9735 17629
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 11348 17669 11376 17700
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12434 17688 12440 17740
rect 12492 17688 12498 17740
rect 13630 17688 13636 17740
rect 13688 17688 13694 17740
rect 14550 17688 14556 17740
rect 14608 17688 14614 17740
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 15470 17728 15476 17740
rect 14792 17700 15476 17728
rect 14792 17688 14798 17700
rect 15470 17688 15476 17700
rect 15528 17688 15534 17740
rect 15654 17688 15660 17740
rect 15712 17688 15718 17740
rect 16132 17737 16160 17768
rect 16316 17768 16856 17796
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 10152 17632 10977 17660
rect 5712 17595 5770 17601
rect 5712 17561 5724 17595
rect 5758 17592 5770 17595
rect 5902 17592 5908 17604
rect 5758 17564 5908 17592
rect 5758 17561 5770 17564
rect 5712 17555 5770 17561
rect 5902 17552 5908 17564
rect 5960 17552 5966 17604
rect 6546 17552 6552 17604
rect 6604 17592 6610 17604
rect 7162 17595 7220 17601
rect 7162 17592 7174 17595
rect 6604 17564 7174 17592
rect 6604 17552 6610 17564
rect 7162 17561 7174 17564
rect 7208 17561 7220 17595
rect 7162 17555 7220 17561
rect 10152 17536 10180 17632
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 10980 17592 11008 17623
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11664 17632 11713 17660
rect 11664 17620 11670 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 12158 17620 12164 17672
rect 12216 17620 12222 17672
rect 15672 17660 15700 17688
rect 16316 17669 16344 17768
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 16758 17688 16764 17740
rect 16816 17688 16822 17740
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 17773 17731 17831 17737
rect 17773 17728 17785 17731
rect 17552 17700 17785 17728
rect 17552 17688 17558 17700
rect 17773 17697 17785 17700
rect 17819 17697 17831 17731
rect 17773 17691 17831 17697
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15672 17632 15853 17660
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16623 17663 16681 17669
rect 16623 17660 16635 17663
rect 16301 17623 16359 17629
rect 16408 17632 16635 17660
rect 11425 17595 11483 17601
rect 11425 17592 11437 17595
rect 10980 17564 11437 17592
rect 11425 17561 11437 17564
rect 11471 17561 11483 17595
rect 11425 17555 11483 17561
rect 11517 17595 11575 17601
rect 11517 17561 11529 17595
rect 11563 17592 11575 17595
rect 12682 17595 12740 17601
rect 12682 17592 12694 17595
rect 11563 17564 11652 17592
rect 11563 17561 11575 17564
rect 11517 17555 11575 17561
rect 11624 17536 11652 17564
rect 12360 17564 12694 17592
rect 6825 17527 6883 17533
rect 6825 17493 6837 17527
rect 6871 17524 6883 17527
rect 8110 17524 8116 17536
rect 6871 17496 8116 17524
rect 6871 17493 6883 17496
rect 6825 17487 6883 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 8294 17484 8300 17536
rect 8352 17484 8358 17536
rect 10134 17484 10140 17536
rect 10192 17484 10198 17536
rect 10410 17484 10416 17536
rect 10468 17484 10474 17536
rect 11149 17527 11207 17533
rect 11149 17493 11161 17527
rect 11195 17524 11207 17527
rect 11330 17524 11336 17536
rect 11195 17496 11336 17524
rect 11195 17493 11207 17496
rect 11149 17487 11207 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11606 17484 11612 17536
rect 11664 17484 11670 17536
rect 12360 17533 12388 17564
rect 12682 17561 12694 17564
rect 12728 17561 12740 17595
rect 12682 17555 12740 17561
rect 14090 17552 14096 17604
rect 14148 17592 14154 17604
rect 14148 17564 15516 17592
rect 14148 17552 14154 17564
rect 12345 17527 12403 17533
rect 12345 17493 12357 17527
rect 12391 17493 12403 17527
rect 12345 17487 12403 17493
rect 13817 17527 13875 17533
rect 13817 17493 13829 17527
rect 13863 17524 13875 17527
rect 14366 17524 14372 17536
rect 13863 17496 14372 17524
rect 13863 17493 13875 17496
rect 13817 17487 13875 17493
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 14458 17484 14464 17536
rect 14516 17484 14522 17536
rect 15488 17524 15516 17564
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 15657 17595 15715 17601
rect 15657 17592 15669 17595
rect 15620 17564 15669 17592
rect 15620 17552 15626 17564
rect 15657 17561 15669 17564
rect 15703 17592 15715 17595
rect 15746 17592 15752 17604
rect 15703 17564 15752 17592
rect 15703 17561 15715 17564
rect 15657 17555 15715 17561
rect 15746 17552 15752 17564
rect 15804 17552 15810 17604
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 16408 17592 16436 17632
rect 16623 17629 16635 17632
rect 16669 17629 16681 17663
rect 16623 17623 16681 17629
rect 17954 17620 17960 17672
rect 18012 17620 18018 17672
rect 18524 17669 18552 17836
rect 18877 17833 18889 17836
rect 18923 17864 18935 17867
rect 19242 17864 19248 17876
rect 18923 17836 19248 17864
rect 18923 17833 18935 17836
rect 18877 17827 18935 17833
rect 19242 17824 19248 17836
rect 19300 17864 19306 17876
rect 19337 17867 19395 17873
rect 19337 17864 19349 17867
rect 19300 17836 19349 17864
rect 19300 17824 19306 17836
rect 19337 17833 19349 17836
rect 19383 17833 19395 17867
rect 19337 17827 19395 17833
rect 19886 17824 19892 17876
rect 19944 17864 19950 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 19944 17836 22569 17864
rect 19944 17824 19950 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 23937 17867 23995 17873
rect 23937 17833 23949 17867
rect 23983 17864 23995 17867
rect 25130 17864 25136 17876
rect 23983 17836 25136 17864
rect 23983 17833 23995 17836
rect 23937 17827 23995 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 26326 17824 26332 17876
rect 26384 17864 26390 17876
rect 27801 17867 27859 17873
rect 27801 17864 27813 17867
rect 26384 17836 27813 17864
rect 26384 17824 26390 17836
rect 27801 17833 27813 17836
rect 27847 17833 27859 17867
rect 27801 17827 27859 17833
rect 18690 17688 18696 17740
rect 18748 17688 18754 17740
rect 18969 17731 19027 17737
rect 18969 17697 18981 17731
rect 19015 17728 19027 17731
rect 19334 17728 19340 17740
rect 19015 17700 19196 17728
rect 19015 17697 19027 17700
rect 18969 17691 19027 17697
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 15988 17564 16436 17592
rect 17313 17595 17371 17601
rect 15988 17552 15994 17564
rect 17313 17561 17325 17595
rect 17359 17592 17371 17595
rect 18230 17592 18236 17604
rect 17359 17564 18236 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 17328 17524 17356 17555
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 18708 17592 18736 17688
rect 19168 17672 19196 17700
rect 19306 17688 19340 17728
rect 19392 17688 19398 17740
rect 19904 17728 19932 17824
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17765 20039 17799
rect 19981 17759 20039 17765
rect 20625 17799 20683 17805
rect 20625 17765 20637 17799
rect 20671 17796 20683 17799
rect 20671 17768 23520 17796
rect 20671 17765 20683 17768
rect 20625 17759 20683 17765
rect 19628 17700 19932 17728
rect 19996 17728 20024 17759
rect 19996 17700 20668 17728
rect 19058 17620 19064 17672
rect 19116 17620 19122 17672
rect 19150 17620 19156 17672
rect 19208 17620 19214 17672
rect 19306 17592 19334 17688
rect 19537 17673 19595 17679
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 19537 17639 19549 17673
rect 19583 17670 19595 17673
rect 19628 17670 19656 17700
rect 19886 17670 19892 17672
rect 19583 17642 19656 17670
rect 19812 17669 19892 17670
rect 19797 17663 19892 17669
rect 19583 17639 19595 17642
rect 19537 17633 19595 17639
rect 19797 17629 19809 17663
rect 19843 17642 19892 17663
rect 19843 17629 19855 17642
rect 19797 17623 19855 17629
rect 19886 17620 19892 17642
rect 19944 17620 19950 17672
rect 20070 17620 20076 17672
rect 20128 17620 20134 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 20180 17632 20361 17660
rect 20180 17592 20208 17632
rect 20349 17629 20361 17632
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17656 20499 17663
rect 20640 17656 20668 17700
rect 21192 17700 21864 17728
rect 21192 17669 21220 17700
rect 21836 17672 21864 17700
rect 23382 17688 23388 17740
rect 23440 17688 23446 17740
rect 23492 17737 23520 17768
rect 23477 17731 23535 17737
rect 23477 17697 23489 17731
rect 23523 17697 23535 17731
rect 23477 17691 23535 17697
rect 25038 17688 25044 17740
rect 25096 17728 25102 17740
rect 26053 17731 26111 17737
rect 26053 17728 26065 17731
rect 25096 17700 26065 17728
rect 25096 17688 25102 17700
rect 26053 17697 26065 17700
rect 26099 17697 26111 17731
rect 26053 17691 26111 17697
rect 20487 17629 20668 17656
rect 20441 17628 20668 17629
rect 21177 17663 21235 17669
rect 21177 17629 21189 17663
rect 21223 17629 21235 17663
rect 20441 17623 20499 17628
rect 21177 17623 21235 17629
rect 21358 17620 21364 17672
rect 21416 17620 21422 17672
rect 21818 17620 21824 17672
rect 21876 17660 21882 17672
rect 21913 17663 21971 17669
rect 21913 17660 21925 17663
rect 21876 17632 21925 17660
rect 21876 17620 21882 17632
rect 21913 17629 21925 17632
rect 21959 17629 21971 17663
rect 21913 17623 21971 17629
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22189 17663 22247 17669
rect 22189 17660 22201 17663
rect 22152 17632 22201 17660
rect 22152 17620 22158 17632
rect 22189 17629 22201 17632
rect 22235 17629 22247 17663
rect 24762 17660 24768 17672
rect 22189 17623 22247 17629
rect 22848 17632 24768 17660
rect 18708 17564 19334 17592
rect 19516 17564 20208 17592
rect 15488 17496 17356 17524
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 17920 17496 18705 17524
rect 17920 17484 17926 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 19516 17524 19544 17564
rect 20254 17552 20260 17604
rect 20312 17552 20318 17604
rect 21726 17552 21732 17604
rect 21784 17552 21790 17604
rect 22278 17552 22284 17604
rect 22336 17592 22342 17604
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22336 17564 22753 17592
rect 22336 17552 22342 17564
rect 22741 17561 22753 17564
rect 22787 17592 22799 17595
rect 22848 17592 22876 17632
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25498 17620 25504 17672
rect 25556 17620 25562 17672
rect 22787 17564 22876 17592
rect 22925 17595 22983 17601
rect 22787 17561 22799 17564
rect 22741 17555 22799 17561
rect 22925 17561 22937 17595
rect 22971 17592 22983 17595
rect 23106 17592 23112 17604
rect 22971 17564 23112 17592
rect 22971 17561 22983 17564
rect 22925 17555 22983 17561
rect 19024 17496 19544 17524
rect 19024 17484 19030 17496
rect 19610 17484 19616 17536
rect 19668 17484 19674 17536
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21361 17527 21419 17533
rect 21361 17524 21373 17527
rect 21140 17496 21373 17524
rect 21140 17484 21146 17496
rect 21361 17493 21373 17496
rect 21407 17493 21419 17527
rect 21361 17487 21419 17493
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 22940 17524 22968 17555
rect 23106 17552 23112 17564
rect 23164 17552 23170 17604
rect 23566 17552 23572 17604
rect 23624 17552 23630 17604
rect 26329 17595 26387 17601
rect 26329 17592 26341 17595
rect 25700 17564 26341 17592
rect 25700 17533 25728 17564
rect 26329 17561 26341 17564
rect 26375 17561 26387 17595
rect 26329 17555 26387 17561
rect 27062 17552 27068 17604
rect 27120 17552 27126 17604
rect 22612 17496 22968 17524
rect 25685 17527 25743 17533
rect 22612 17484 22618 17496
rect 25685 17493 25697 17527
rect 25731 17493 25743 17527
rect 25685 17487 25743 17493
rect 1104 17434 31280 17456
rect 1104 17382 4922 17434
rect 4974 17382 4986 17434
rect 5038 17382 5050 17434
rect 5102 17382 5114 17434
rect 5166 17382 5178 17434
rect 5230 17382 5242 17434
rect 5294 17382 10922 17434
rect 10974 17382 10986 17434
rect 11038 17382 11050 17434
rect 11102 17382 11114 17434
rect 11166 17382 11178 17434
rect 11230 17382 11242 17434
rect 11294 17382 16922 17434
rect 16974 17382 16986 17434
rect 17038 17382 17050 17434
rect 17102 17382 17114 17434
rect 17166 17382 17178 17434
rect 17230 17382 17242 17434
rect 17294 17382 22922 17434
rect 22974 17382 22986 17434
rect 23038 17382 23050 17434
rect 23102 17382 23114 17434
rect 23166 17382 23178 17434
rect 23230 17382 23242 17434
rect 23294 17382 28922 17434
rect 28974 17382 28986 17434
rect 29038 17382 29050 17434
rect 29102 17382 29114 17434
rect 29166 17382 29178 17434
rect 29230 17382 29242 17434
rect 29294 17382 31280 17434
rect 1104 17360 31280 17382
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6546 17320 6552 17332
rect 5951 17292 6552 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6788 17292 6837 17320
rect 6788 17280 6794 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 8294 17320 8300 17332
rect 6825 17283 6883 17289
rect 7852 17292 8300 17320
rect 7852 17252 7880 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8444 17292 10088 17320
rect 8444 17280 8450 17292
rect 7852 17224 8064 17252
rect 7852 17193 7880 17224
rect 8036 17193 8064 17224
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 9024 17255 9082 17261
rect 8168 17224 8340 17252
rect 8168 17212 8174 17224
rect 5721 17187 5779 17193
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 6733 17187 6791 17193
rect 5767 17156 6408 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 6380 17057 6408 17156
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6779 17156 7205 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7193 17153 7205 17156
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 8022 17187 8080 17193
rect 8022 17153 8034 17187
rect 8068 17153 8080 17187
rect 8022 17147 8080 17153
rect 6454 17076 6460 17128
rect 6512 17076 6518 17128
rect 6822 17076 6828 17128
rect 6880 17116 6886 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6880 17088 6929 17116
rect 6880 17076 6886 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 6365 17051 6423 17057
rect 6365 17017 6377 17051
rect 6411 17017 6423 17051
rect 6472 17048 6500 17076
rect 7944 17048 7972 17147
rect 8202 17144 8208 17196
rect 8260 17144 8266 17196
rect 8312 17193 8340 17224
rect 8680 17224 8892 17252
rect 8478 17193 8484 17196
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8435 17187 8484 17193
rect 8435 17153 8447 17187
rect 8481 17153 8484 17187
rect 8435 17147 8484 17153
rect 8478 17144 8484 17147
rect 8536 17184 8542 17196
rect 8680 17184 8708 17224
rect 8536 17156 8708 17184
rect 8536 17144 8542 17156
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 8864 17184 8892 17224
rect 9024 17221 9036 17255
rect 9070 17252 9082 17255
rect 9122 17252 9128 17264
rect 9070 17224 9128 17252
rect 9070 17221 9082 17224
rect 9024 17215 9082 17221
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 9582 17212 9588 17264
rect 9640 17252 9646 17264
rect 10060 17252 10088 17292
rect 10134 17280 10140 17332
rect 10192 17280 10198 17332
rect 10410 17280 10416 17332
rect 10468 17320 10474 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 10468 17292 10701 17320
rect 10468 17280 10474 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 11664 17292 11744 17320
rect 11664 17280 11670 17292
rect 9640 17224 9987 17252
rect 10060 17224 10548 17252
rect 9640 17212 9646 17224
rect 9959 17184 9987 17224
rect 10520 17184 10548 17224
rect 10594 17212 10600 17264
rect 10652 17212 10658 17264
rect 11716 17252 11744 17292
rect 12158 17280 12164 17332
rect 12216 17320 12222 17332
rect 12989 17323 13047 17329
rect 12989 17320 13001 17323
rect 12216 17292 13001 17320
rect 12216 17280 12222 17292
rect 12989 17289 13001 17292
rect 13035 17289 13047 17323
rect 12989 17283 13047 17289
rect 15194 17280 15200 17332
rect 15252 17280 15258 17332
rect 16666 17280 16672 17332
rect 16724 17320 16730 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16724 17292 17141 17320
rect 16724 17280 16730 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 17129 17283 17187 17289
rect 18414 17280 18420 17332
rect 18472 17280 18478 17332
rect 19518 17280 19524 17332
rect 19576 17280 19582 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 20809 17323 20867 17329
rect 20809 17320 20821 17323
rect 20312 17292 20821 17320
rect 20312 17280 20318 17292
rect 20809 17289 20821 17292
rect 20855 17289 20867 17323
rect 23385 17323 23443 17329
rect 23385 17320 23397 17323
rect 20809 17283 20867 17289
rect 20916 17292 23397 17320
rect 15102 17252 15108 17264
rect 11716 17224 15108 17252
rect 15102 17212 15108 17224
rect 15160 17212 15166 17264
rect 16758 17212 16764 17264
rect 16816 17252 16822 17264
rect 17037 17255 17095 17261
rect 17037 17252 17049 17255
rect 16816 17224 17049 17252
rect 16816 17212 16822 17224
rect 17037 17221 17049 17224
rect 17083 17221 17095 17255
rect 17037 17215 17095 17221
rect 17678 17212 17684 17264
rect 17736 17212 17742 17264
rect 19058 17212 19064 17264
rect 19116 17252 19122 17264
rect 20916 17252 20944 17292
rect 23385 17289 23397 17292
rect 23431 17289 23443 17323
rect 23385 17283 23443 17289
rect 24026 17280 24032 17332
rect 24084 17280 24090 17332
rect 24397 17323 24455 17329
rect 24397 17289 24409 17323
rect 24443 17289 24455 17323
rect 24397 17283 24455 17289
rect 19116 17224 20944 17252
rect 19116 17212 19122 17224
rect 21358 17212 21364 17264
rect 21416 17252 21422 17264
rect 21821 17255 21879 17261
rect 21821 17252 21833 17255
rect 21416 17224 21833 17252
rect 21416 17212 21422 17224
rect 21821 17221 21833 17224
rect 21867 17221 21879 17255
rect 21821 17215 21879 17221
rect 22646 17212 22652 17264
rect 22704 17252 22710 17264
rect 23474 17252 23480 17264
rect 22704 17224 23480 17252
rect 22704 17212 22710 17224
rect 23474 17212 23480 17224
rect 23532 17212 23538 17264
rect 24044 17252 24072 17280
rect 23584 17224 24072 17252
rect 24412 17252 24440 17283
rect 24762 17280 24768 17332
rect 24820 17320 24826 17332
rect 24857 17323 24915 17329
rect 24857 17320 24869 17323
rect 24820 17292 24869 17320
rect 24820 17280 24826 17292
rect 24857 17289 24869 17292
rect 24903 17289 24915 17323
rect 24857 17283 24915 17289
rect 25225 17323 25283 17329
rect 25225 17289 25237 17323
rect 25271 17320 25283 17323
rect 25498 17320 25504 17332
rect 25271 17292 25504 17320
rect 25271 17289 25283 17292
rect 25225 17283 25283 17289
rect 25498 17280 25504 17292
rect 25556 17280 25562 17332
rect 24412 17224 25360 17252
rect 11422 17184 11428 17196
rect 8864 17156 9812 17184
rect 9959 17156 10364 17184
rect 10520 17156 11428 17184
rect 9784 17116 9812 17156
rect 10042 17116 10048 17128
rect 9784 17088 10048 17116
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 6472 17020 7972 17048
rect 10229 17051 10287 17057
rect 6365 17011 6423 17017
rect 10229 17017 10241 17051
rect 10275 17048 10287 17051
rect 10336 17048 10364 17156
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 11514 17144 11520 17196
rect 11572 17144 11578 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17184 13415 17187
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13403 17156 13829 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11716 17116 11744 17147
rect 14366 17144 14372 17196
rect 14424 17144 14430 17196
rect 16482 17144 16488 17196
rect 16540 17144 16546 17196
rect 17862 17184 17868 17196
rect 17236 17156 17868 17184
rect 11204 17088 11744 17116
rect 11204 17076 11210 17088
rect 13446 17076 13452 17128
rect 13504 17076 13510 17128
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 13688 17088 15148 17116
rect 13688 17076 13694 17088
rect 10275 17020 10364 17048
rect 15120 17048 15148 17088
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17236 17125 17264 17156
rect 17862 17144 17868 17156
rect 17920 17184 17926 17196
rect 17957 17187 18015 17193
rect 17957 17184 17969 17187
rect 17920 17156 17969 17184
rect 17920 17144 17926 17156
rect 17957 17153 17969 17156
rect 18003 17153 18015 17187
rect 17957 17147 18015 17153
rect 18138 17144 18144 17196
rect 18196 17190 18202 17196
rect 18233 17190 18291 17193
rect 18196 17187 18291 17190
rect 18196 17162 18245 17187
rect 18196 17144 18202 17162
rect 18233 17153 18245 17162
rect 18279 17153 18291 17187
rect 18509 17187 18567 17193
rect 18509 17184 18521 17187
rect 18233 17147 18291 17153
rect 18432 17156 18521 17184
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 16632 17088 17233 17116
rect 16632 17076 16638 17088
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17402 17048 17408 17060
rect 15120 17020 17408 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 18248 17048 18276 17147
rect 18432 17128 18460 17156
rect 18509 17153 18521 17156
rect 18555 17153 18567 17187
rect 19153 17187 19211 17193
rect 19153 17184 19165 17187
rect 18509 17147 18567 17153
rect 18984 17156 19165 17184
rect 18984 17128 19012 17156
rect 19153 17153 19165 17156
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 19242 17144 19248 17196
rect 19300 17144 19306 17196
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17184 21051 17187
rect 22094 17184 22100 17196
rect 21039 17156 22100 17184
rect 21039 17153 21051 17156
rect 20993 17147 21051 17153
rect 22094 17144 22100 17156
rect 22152 17144 22158 17196
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 22922 17184 22928 17196
rect 22612 17156 22928 17184
rect 22612 17144 22618 17156
rect 22922 17144 22928 17156
rect 22980 17144 22986 17196
rect 23584 17193 23612 17224
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17153 23627 17187
rect 23569 17147 23627 17153
rect 23658 17144 23664 17196
rect 23716 17184 23722 17196
rect 25332 17193 25360 17224
rect 24029 17187 24087 17193
rect 24029 17184 24041 17187
rect 23716 17156 24041 17184
rect 23716 17144 23722 17156
rect 24029 17153 24041 17156
rect 24075 17153 24087 17187
rect 24029 17147 24087 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17153 25375 17187
rect 25317 17147 25375 17153
rect 26970 17144 26976 17196
rect 27028 17184 27034 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 27028 17156 27169 17184
rect 27028 17144 27034 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 18414 17076 18420 17128
rect 18472 17076 18478 17128
rect 18966 17076 18972 17128
rect 19024 17076 19030 17128
rect 19058 17076 19064 17128
rect 19116 17076 19122 17128
rect 19337 17119 19395 17125
rect 19337 17085 19349 17119
rect 19383 17085 19395 17119
rect 19337 17079 19395 17085
rect 19352 17048 19380 17079
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 20956 17088 21097 17116
rect 20956 17076 20962 17088
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 21085 17079 21143 17085
rect 21177 17119 21235 17125
rect 21177 17085 21189 17119
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 17972 17020 18184 17048
rect 18248 17020 19380 17048
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 8619 16952 11529 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 11517 16943 11575 16949
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 12250 16980 12256 16992
rect 11931 16952 12256 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 16758 16940 16764 16992
rect 16816 16980 16822 16992
rect 17972 16980 18000 17020
rect 16816 16952 18000 16980
rect 16816 16940 16822 16952
rect 18046 16940 18052 16992
rect 18104 16940 18110 16992
rect 18156 16980 18184 17020
rect 20714 16980 20720 16992
rect 18156 16952 20720 16980
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 20916 16980 20944 17076
rect 20990 17008 20996 17060
rect 21048 17048 21054 17060
rect 21192 17048 21220 17079
rect 21266 17076 21272 17128
rect 21324 17116 21330 17128
rect 22189 17119 22247 17125
rect 22189 17116 22201 17119
rect 21324 17088 22201 17116
rect 21324 17076 21330 17088
rect 22189 17085 22201 17088
rect 22235 17116 22247 17119
rect 22235 17088 22416 17116
rect 22235 17085 22247 17088
rect 22189 17079 22247 17085
rect 22097 17051 22155 17057
rect 22097 17048 22109 17051
rect 21048 17020 22109 17048
rect 21048 17008 21054 17020
rect 22097 17017 22109 17020
rect 22143 17048 22155 17051
rect 22278 17048 22284 17060
rect 22143 17020 22284 17048
rect 22143 17017 22155 17020
rect 22097 17011 22155 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22388 17048 22416 17088
rect 23014 17076 23020 17128
rect 23072 17116 23078 17128
rect 23382 17116 23388 17128
rect 23072 17088 23388 17116
rect 23072 17076 23078 17088
rect 23382 17076 23388 17088
rect 23440 17116 23446 17128
rect 23753 17119 23811 17125
rect 23753 17116 23765 17119
rect 23440 17088 23765 17116
rect 23440 17076 23446 17088
rect 23753 17085 23765 17088
rect 23799 17085 23811 17119
rect 23753 17079 23811 17085
rect 23566 17048 23572 17060
rect 22388 17020 23572 17048
rect 23566 17008 23572 17020
rect 23624 17008 23630 17060
rect 23768 17048 23796 17079
rect 23934 17076 23940 17128
rect 23992 17076 23998 17128
rect 24581 17119 24639 17125
rect 24581 17085 24593 17119
rect 24627 17085 24639 17119
rect 24581 17079 24639 17085
rect 24765 17119 24823 17125
rect 24765 17085 24777 17119
rect 24811 17116 24823 17119
rect 24811 17088 24900 17116
rect 24811 17085 24823 17088
rect 24765 17079 24823 17085
rect 24596 17048 24624 17079
rect 24872 17060 24900 17088
rect 23768 17020 24624 17048
rect 24854 17008 24860 17060
rect 24912 17008 24918 17060
rect 22002 16989 22008 16992
rect 21986 16983 22008 16989
rect 21986 16980 21998 16983
rect 20916 16952 21998 16980
rect 21986 16949 21998 16952
rect 21986 16943 22008 16949
rect 22002 16940 22008 16943
rect 22060 16940 22066 16992
rect 22465 16983 22523 16989
rect 22465 16949 22477 16983
rect 22511 16980 22523 16983
rect 22646 16980 22652 16992
rect 22511 16952 22652 16980
rect 22511 16949 22523 16952
rect 22465 16943 22523 16949
rect 22646 16940 22652 16952
rect 22704 16940 22710 16992
rect 25498 16940 25504 16992
rect 25556 16940 25562 16992
rect 27065 16983 27123 16989
rect 27065 16949 27077 16983
rect 27111 16980 27123 16983
rect 27154 16980 27160 16992
rect 27111 16952 27160 16980
rect 27111 16949 27123 16952
rect 27065 16943 27123 16949
rect 27154 16940 27160 16952
rect 27212 16940 27218 16992
rect 1104 16890 31280 16912
rect 1104 16838 4182 16890
rect 4234 16838 4246 16890
rect 4298 16838 4310 16890
rect 4362 16838 4374 16890
rect 4426 16838 4438 16890
rect 4490 16838 4502 16890
rect 4554 16838 10182 16890
rect 10234 16838 10246 16890
rect 10298 16838 10310 16890
rect 10362 16838 10374 16890
rect 10426 16838 10438 16890
rect 10490 16838 10502 16890
rect 10554 16838 16182 16890
rect 16234 16838 16246 16890
rect 16298 16838 16310 16890
rect 16362 16838 16374 16890
rect 16426 16838 16438 16890
rect 16490 16838 16502 16890
rect 16554 16838 22182 16890
rect 22234 16838 22246 16890
rect 22298 16838 22310 16890
rect 22362 16838 22374 16890
rect 22426 16838 22438 16890
rect 22490 16838 22502 16890
rect 22554 16838 28182 16890
rect 28234 16838 28246 16890
rect 28298 16838 28310 16890
rect 28362 16838 28374 16890
rect 28426 16838 28438 16890
rect 28490 16838 28502 16890
rect 28554 16838 31280 16890
rect 1104 16816 31280 16838
rect 3878 16776 3884 16788
rect 3068 16748 3884 16776
rect 3068 16649 3096 16748
rect 3878 16736 3884 16748
rect 3936 16776 3942 16788
rect 8018 16776 8024 16788
rect 3936 16748 8024 16776
rect 3936 16736 3942 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9122 16736 9128 16788
rect 9180 16736 9186 16788
rect 11146 16736 11152 16788
rect 11204 16736 11210 16788
rect 14090 16776 14096 16788
rect 11440 16748 14096 16776
rect 6822 16668 6828 16720
rect 6880 16708 6886 16720
rect 11440 16708 11468 16748
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14366 16736 14372 16788
rect 14424 16736 14430 16788
rect 15841 16779 15899 16785
rect 15841 16745 15853 16779
rect 15887 16776 15899 16779
rect 15930 16776 15936 16788
rect 15887 16748 15936 16776
rect 15887 16745 15899 16748
rect 15841 16739 15899 16745
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 18046 16736 18052 16788
rect 18104 16736 18110 16788
rect 19058 16736 19064 16788
rect 19116 16736 19122 16788
rect 19426 16736 19432 16788
rect 19484 16736 19490 16788
rect 20714 16736 20720 16788
rect 20772 16776 20778 16788
rect 21726 16776 21732 16788
rect 20772 16748 21732 16776
rect 20772 16736 20778 16748
rect 21726 16736 21732 16748
rect 21784 16736 21790 16788
rect 22370 16736 22376 16788
rect 22428 16776 22434 16788
rect 23014 16776 23020 16788
rect 22428 16748 23020 16776
rect 22428 16736 22434 16748
rect 23014 16736 23020 16748
rect 23072 16736 23078 16788
rect 23106 16736 23112 16788
rect 23164 16776 23170 16788
rect 23661 16779 23719 16785
rect 23164 16748 23520 16776
rect 23164 16736 23170 16748
rect 6880 16680 11468 16708
rect 6880 16668 6886 16680
rect 11514 16668 11520 16720
rect 11572 16708 11578 16720
rect 11572 16680 11928 16708
rect 11572 16668 11578 16680
rect 11900 16652 11928 16680
rect 3053 16643 3111 16649
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 4614 16640 4620 16652
rect 3292 16612 4620 16640
rect 3292 16600 3298 16612
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 11422 16640 11428 16652
rect 10705 16612 11428 16640
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16541 2559 16575
rect 2501 16535 2559 16541
rect 2314 16396 2320 16448
rect 2372 16396 2378 16448
rect 2516 16436 2544 16535
rect 4338 16532 4344 16584
rect 4396 16532 4402 16584
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16572 9367 16575
rect 9600 16572 9628 16600
rect 10705 16581 10733 16612
rect 11422 16600 11428 16612
rect 11480 16640 11486 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11480 16612 11805 16640
rect 11480 16600 11486 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 11940 16612 14044 16640
rect 11940 16600 11946 16612
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 9355 16544 9628 16572
rect 10428 16544 10517 16572
rect 9355 16541 9367 16544
rect 9309 16535 9367 16541
rect 2961 16507 3019 16513
rect 2961 16473 2973 16507
rect 3007 16504 3019 16507
rect 3789 16507 3847 16513
rect 3789 16504 3801 16507
rect 3007 16476 3801 16504
rect 3007 16473 3019 16476
rect 2961 16467 3019 16473
rect 3789 16473 3801 16476
rect 3835 16473 3847 16507
rect 3789 16467 3847 16473
rect 2593 16439 2651 16445
rect 2593 16436 2605 16439
rect 2516 16408 2605 16436
rect 2593 16405 2605 16408
rect 2639 16405 2651 16439
rect 10428 16436 10456 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 10653 16575 10733 16581
rect 10653 16541 10665 16575
rect 10699 16544 10733 16575
rect 11011 16575 11069 16581
rect 10699 16541 10711 16544
rect 10653 16535 10711 16541
rect 11011 16541 11023 16575
rect 11057 16572 11069 16575
rect 11698 16572 11704 16584
rect 11057 16544 11704 16572
rect 11057 16541 11069 16544
rect 11011 16535 11069 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 10778 16464 10784 16516
rect 10836 16464 10842 16516
rect 10873 16507 10931 16513
rect 10873 16473 10885 16507
rect 10919 16504 10931 16507
rect 10919 16476 11928 16504
rect 10919 16473 10931 16476
rect 10873 16467 10931 16473
rect 11900 16448 11928 16476
rect 11146 16436 11152 16448
rect 10428 16408 11152 16436
rect 2593 16399 2651 16405
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 11241 16439 11299 16445
rect 11241 16405 11253 16439
rect 11287 16436 11299 16439
rect 11330 16436 11336 16448
rect 11287 16408 11336 16436
rect 11287 16405 11299 16408
rect 11241 16399 11299 16405
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 11882 16396 11888 16448
rect 11940 16396 11946 16448
rect 14016 16436 14044 16612
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14384 16572 14412 16736
rect 15286 16640 15292 16652
rect 14476 16612 15292 16640
rect 14476 16581 14504 16612
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 16040 16612 16620 16640
rect 16040 16584 16068 16612
rect 14139 16544 14412 16572
rect 14461 16575 14519 16581
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14461 16541 14473 16575
rect 14507 16541 14519 16575
rect 14461 16535 14519 16541
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 14277 16507 14335 16513
rect 14277 16504 14289 16507
rect 14240 16476 14289 16504
rect 14240 16464 14246 16476
rect 14277 16473 14289 16476
rect 14323 16473 14335 16507
rect 14277 16467 14335 16473
rect 14366 16464 14372 16516
rect 14424 16464 14430 16516
rect 14476 16436 14504 16535
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 14792 16544 15976 16572
rect 14792 16532 14798 16544
rect 15473 16507 15531 16513
rect 15473 16473 15485 16507
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 14016 16408 14504 16436
rect 14645 16439 14703 16445
rect 14645 16405 14657 16439
rect 14691 16436 14703 16439
rect 15194 16436 15200 16448
rect 14691 16408 15200 16436
rect 14691 16405 14703 16408
rect 14645 16399 14703 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15488 16436 15516 16467
rect 15654 16464 15660 16516
rect 15712 16464 15718 16516
rect 15948 16504 15976 16544
rect 16022 16532 16028 16584
rect 16080 16532 16086 16584
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16541 16359 16575
rect 16301 16535 16359 16541
rect 16316 16504 16344 16535
rect 15948 16476 16344 16504
rect 16592 16504 16620 16612
rect 16684 16581 16712 16736
rect 17405 16711 17463 16717
rect 17405 16677 17417 16711
rect 17451 16708 17463 16711
rect 17586 16708 17592 16720
rect 17451 16680 17592 16708
rect 17451 16677 17463 16680
rect 17405 16671 17463 16677
rect 17586 16668 17592 16680
rect 17644 16668 17650 16720
rect 18064 16640 18092 16736
rect 19076 16708 19104 16736
rect 19613 16711 19671 16717
rect 19613 16708 19625 16711
rect 19076 16680 19625 16708
rect 19613 16677 19625 16680
rect 19659 16677 19671 16711
rect 19613 16671 19671 16677
rect 22741 16711 22799 16717
rect 22741 16677 22753 16711
rect 22787 16708 22799 16711
rect 23198 16708 23204 16720
rect 22787 16680 23204 16708
rect 22787 16677 22799 16680
rect 22741 16671 22799 16677
rect 18414 16640 18420 16652
rect 17512 16612 18092 16640
rect 18156 16612 18420 16640
rect 17512 16581 17540 16612
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 16776 16504 16804 16535
rect 16592 16476 16804 16504
rect 15746 16436 15752 16448
rect 15488 16408 15752 16436
rect 15746 16396 15752 16408
rect 15804 16436 15810 16448
rect 18156 16436 18184 16612
rect 18414 16600 18420 16612
rect 18472 16600 18478 16652
rect 19242 16640 19248 16652
rect 18800 16612 19248 16640
rect 18690 16532 18696 16584
rect 18748 16532 18754 16584
rect 18800 16581 18828 16612
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19628 16640 19656 16671
rect 23198 16668 23204 16680
rect 23256 16668 23262 16720
rect 23492 16708 23520 16748
rect 23661 16745 23673 16779
rect 23707 16776 23719 16779
rect 23934 16776 23940 16788
rect 23707 16748 23940 16776
rect 23707 16745 23719 16748
rect 23661 16739 23719 16745
rect 23934 16736 23940 16748
rect 23992 16736 23998 16788
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 26126 16779 26184 16785
rect 26126 16776 26138 16779
rect 25556 16748 26138 16776
rect 25556 16736 25562 16748
rect 26126 16745 26138 16748
rect 26172 16745 26184 16779
rect 26126 16739 26184 16745
rect 27614 16736 27620 16788
rect 27672 16736 27678 16788
rect 23566 16708 23572 16720
rect 23492 16680 23572 16708
rect 23492 16649 23520 16680
rect 23566 16668 23572 16680
rect 23624 16708 23630 16720
rect 23624 16680 24716 16708
rect 23624 16668 23630 16680
rect 23293 16643 23351 16649
rect 23293 16640 23305 16643
rect 19628 16612 20760 16640
rect 20732 16581 20760 16612
rect 20824 16612 23305 16640
rect 18785 16575 18843 16581
rect 18785 16541 18797 16575
rect 18831 16541 18843 16575
rect 18785 16535 18843 16541
rect 18969 16575 19027 16581
rect 18969 16541 18981 16575
rect 19015 16541 19027 16575
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 18969 16535 19027 16541
rect 19168 16544 19717 16572
rect 18708 16504 18736 16532
rect 18984 16504 19012 16535
rect 18708 16476 19012 16504
rect 19168 16448 19196 16544
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 19242 16464 19248 16516
rect 19300 16504 19306 16516
rect 19797 16507 19855 16513
rect 19797 16504 19809 16507
rect 19300 16476 19809 16504
rect 19300 16464 19306 16476
rect 19797 16473 19809 16476
rect 19843 16504 19855 16507
rect 20070 16504 20076 16516
rect 19843 16476 20076 16504
rect 19843 16473 19855 16476
rect 19797 16467 19855 16473
rect 20070 16464 20076 16476
rect 20128 16504 20134 16516
rect 20824 16504 20852 16612
rect 23293 16609 23305 16612
rect 23339 16609 23351 16643
rect 23293 16603 23351 16609
rect 23477 16643 23535 16649
rect 23477 16609 23489 16643
rect 23523 16609 23535 16643
rect 23477 16603 23535 16609
rect 24394 16600 24400 16652
rect 24452 16600 24458 16652
rect 24688 16649 24716 16680
rect 24673 16643 24731 16649
rect 24673 16609 24685 16643
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16640 25927 16643
rect 26234 16640 26240 16652
rect 25915 16612 26240 16640
rect 25915 16609 25927 16612
rect 25869 16603 25927 16609
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 20901 16575 20959 16581
rect 20901 16541 20913 16575
rect 20947 16572 20959 16575
rect 22094 16572 22100 16584
rect 20947 16544 22100 16572
rect 20947 16541 20959 16544
rect 20901 16535 20959 16541
rect 22094 16532 22100 16544
rect 22152 16532 22158 16584
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23106 16572 23112 16584
rect 23063 16544 23112 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23198 16532 23204 16584
rect 23256 16532 23262 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23845 16575 23903 16581
rect 23845 16541 23857 16575
rect 23891 16572 23903 16575
rect 24026 16572 24032 16584
rect 23891 16544 24032 16572
rect 23891 16541 23903 16544
rect 23845 16535 23903 16541
rect 21358 16504 21364 16516
rect 20128 16476 20852 16504
rect 20916 16476 21364 16504
rect 20128 16464 20134 16476
rect 15804 16408 18184 16436
rect 15804 16396 15810 16408
rect 18782 16396 18788 16448
rect 18840 16396 18846 16448
rect 19150 16396 19156 16448
rect 19208 16396 19214 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 19445 16439 19503 16445
rect 19445 16436 19457 16439
rect 19392 16408 19457 16436
rect 19392 16396 19398 16408
rect 19445 16405 19457 16408
rect 19491 16436 19503 16439
rect 19886 16436 19892 16448
rect 19491 16408 19892 16436
rect 19491 16405 19503 16408
rect 19445 16399 19503 16405
rect 19886 16396 19892 16408
rect 19944 16396 19950 16448
rect 20809 16439 20867 16445
rect 20809 16405 20821 16439
rect 20855 16436 20867 16439
rect 20916 16436 20944 16476
rect 21358 16464 21364 16476
rect 21416 16464 21422 16516
rect 22741 16507 22799 16513
rect 22741 16473 22753 16507
rect 22787 16473 22799 16507
rect 22940 16504 22968 16532
rect 23400 16504 23428 16535
rect 24026 16532 24032 16544
rect 24084 16532 24090 16584
rect 24762 16532 24768 16584
rect 24820 16532 24826 16584
rect 27154 16532 27160 16584
rect 27212 16572 27218 16584
rect 27212 16544 27278 16572
rect 27212 16532 27218 16544
rect 22940 16476 23428 16504
rect 24213 16507 24271 16513
rect 22741 16467 22799 16473
rect 24213 16473 24225 16507
rect 24259 16504 24271 16507
rect 24302 16504 24308 16516
rect 24259 16476 24308 16504
rect 24259 16473 24271 16476
rect 24213 16467 24271 16473
rect 20855 16408 20944 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 22756 16436 22784 16467
rect 24302 16464 24308 16476
rect 24360 16464 24366 16516
rect 26510 16436 26516 16448
rect 21048 16408 26516 16436
rect 21048 16396 21054 16408
rect 26510 16396 26516 16408
rect 26568 16396 26574 16448
rect 1104 16346 31280 16368
rect 1104 16294 4922 16346
rect 4974 16294 4986 16346
rect 5038 16294 5050 16346
rect 5102 16294 5114 16346
rect 5166 16294 5178 16346
rect 5230 16294 5242 16346
rect 5294 16294 10922 16346
rect 10974 16294 10986 16346
rect 11038 16294 11050 16346
rect 11102 16294 11114 16346
rect 11166 16294 11178 16346
rect 11230 16294 11242 16346
rect 11294 16294 16922 16346
rect 16974 16294 16986 16346
rect 17038 16294 17050 16346
rect 17102 16294 17114 16346
rect 17166 16294 17178 16346
rect 17230 16294 17242 16346
rect 17294 16294 22922 16346
rect 22974 16294 22986 16346
rect 23038 16294 23050 16346
rect 23102 16294 23114 16346
rect 23166 16294 23178 16346
rect 23230 16294 23242 16346
rect 23294 16294 28922 16346
rect 28974 16294 28986 16346
rect 29038 16294 29050 16346
rect 29102 16294 29114 16346
rect 29166 16294 29178 16346
rect 29230 16294 29242 16346
rect 29294 16294 31280 16346
rect 1104 16272 31280 16294
rect 3329 16235 3387 16241
rect 3329 16201 3341 16235
rect 3375 16232 3387 16235
rect 4338 16232 4344 16244
rect 3375 16204 4344 16232
rect 3375 16201 3387 16204
rect 3329 16195 3387 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 6638 16192 6644 16244
rect 6696 16232 6702 16244
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 6696 16204 6837 16232
rect 6696 16192 6702 16204
rect 6825 16201 6837 16204
rect 6871 16232 6883 16235
rect 8386 16232 8392 16244
rect 6871 16204 8392 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8665 16235 8723 16241
rect 8665 16201 8677 16235
rect 8711 16201 8723 16235
rect 8665 16195 8723 16201
rect 10229 16235 10287 16241
rect 10229 16201 10241 16235
rect 10275 16201 10287 16235
rect 10229 16195 10287 16201
rect 2216 16167 2274 16173
rect 2216 16133 2228 16167
rect 2262 16164 2274 16167
rect 2314 16164 2320 16176
rect 2262 16136 2320 16164
rect 2262 16133 2274 16136
rect 2216 16127 2274 16133
rect 2314 16124 2320 16136
rect 2372 16124 2378 16176
rect 3878 16124 3884 16176
rect 3936 16124 3942 16176
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 3789 16099 3847 16105
rect 1719 16068 3464 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1946 15988 1952 16040
rect 2004 15988 2010 16040
rect 3436 15969 3464 16068
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 4249 16099 4307 16105
rect 4249 16096 4261 16099
rect 3835 16068 4261 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4249 16065 4261 16068
rect 4295 16065 4307 16099
rect 4356 16096 4384 16192
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 5169 16167 5227 16173
rect 5169 16164 5181 16167
rect 4764 16136 5181 16164
rect 4764 16124 4770 16136
rect 5169 16133 5181 16136
rect 5215 16133 5227 16167
rect 8680 16164 8708 16195
rect 9002 16167 9060 16173
rect 9002 16164 9014 16167
rect 8680 16136 9014 16164
rect 5169 16127 5227 16133
rect 9002 16133 9014 16136
rect 9048 16133 9060 16167
rect 9002 16127 9060 16133
rect 4985 16099 5043 16105
rect 4985 16096 4997 16099
rect 4356 16068 4997 16096
rect 4249 16059 4307 16065
rect 4985 16065 4997 16068
rect 5031 16065 5043 16099
rect 4985 16059 5043 16065
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 5442 16096 5448 16108
rect 5399 16068 5448 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 3970 15988 3976 16040
rect 4028 15988 4034 16040
rect 4801 16031 4859 16037
rect 4801 15997 4813 16031
rect 4847 16028 4859 16031
rect 5276 16028 5304 16059
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6779 16068 7205 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 10244 16096 10272 16195
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10376 16204 10609 16232
rect 10376 16192 10382 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 10689 16235 10747 16241
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 11330 16232 11336 16244
rect 10735 16204 11336 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 10612 16164 10640 16195
rect 11330 16192 11336 16204
rect 11388 16192 11394 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 16758 16232 16764 16244
rect 15712 16204 16764 16232
rect 15712 16192 15718 16204
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 18138 16192 18144 16244
rect 18196 16232 18202 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 18196 16204 18245 16232
rect 18196 16192 18202 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 18233 16195 18291 16201
rect 10962 16164 10968 16176
rect 10612 16136 10968 16164
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 16022 16164 16028 16176
rect 13004 16136 16028 16164
rect 11977 16099 12035 16105
rect 8527 16068 10272 16096
rect 10796 16068 11928 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 4847 16000 5304 16028
rect 4847 15997 4859 16000
rect 4801 15991 4859 15997
rect 3421 15963 3479 15969
rect 3421 15929 3433 15963
rect 3467 15929 3479 15963
rect 3421 15923 3479 15929
rect 1854 15852 1860 15904
rect 1912 15852 1918 15904
rect 3234 15852 3240 15904
rect 3292 15892 3298 15904
rect 3988 15892 4016 15988
rect 4816 15904 4844 15991
rect 6822 15988 6828 16040
rect 6880 16028 6886 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6880 16000 6929 16028
rect 6880 15988 6886 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 7834 15988 7840 16040
rect 7892 15988 7898 16040
rect 7926 15988 7932 16040
rect 7984 16028 7990 16040
rect 8757 16031 8815 16037
rect 8757 16028 8769 16031
rect 7984 16000 8769 16028
rect 7984 15988 7990 16000
rect 8757 15997 8769 16000
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10796 16037 10824 16068
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 9824 16000 10793 16028
rect 9824 15988 9830 16000
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 11422 15988 11428 16040
rect 11480 15988 11486 16040
rect 5537 15963 5595 15969
rect 5537 15929 5549 15963
rect 5583 15960 5595 15963
rect 7282 15960 7288 15972
rect 5583 15932 7288 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 10137 15963 10195 15969
rect 10137 15929 10149 15963
rect 10183 15960 10195 15963
rect 11440 15960 11468 15988
rect 10183 15932 11468 15960
rect 11900 15960 11928 16068
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12618 16096 12624 16108
rect 12023 16068 12624 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13004 16105 13032 16136
rect 16022 16124 16028 16136
rect 16080 16164 16086 16176
rect 18248 16164 18276 16195
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 18506 16232 18512 16244
rect 18380 16204 18512 16232
rect 18380 16192 18386 16204
rect 18506 16192 18512 16204
rect 18564 16232 18570 16244
rect 18564 16204 18736 16232
rect 18564 16192 18570 16204
rect 16080 16136 17724 16164
rect 18248 16136 18644 16164
rect 16080 16124 16086 16136
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 14734 15960 14740 15972
rect 11900 15932 14740 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 14734 15920 14740 15932
rect 14792 15920 14798 15972
rect 3292 15864 4016 15892
rect 3292 15852 3298 15864
rect 4798 15852 4804 15904
rect 4856 15852 4862 15904
rect 6362 15852 6368 15904
rect 6420 15852 6426 15904
rect 12158 15852 12164 15904
rect 12216 15852 12222 15904
rect 12802 15852 12808 15904
rect 12860 15852 12866 15904
rect 13173 15895 13231 15901
rect 13173 15861 13185 15895
rect 13219 15892 13231 15895
rect 14826 15892 14832 15904
rect 13219 15864 14832 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 14826 15852 14832 15864
rect 14884 15892 14890 15904
rect 15102 15892 15108 15904
rect 14884 15864 15108 15892
rect 14884 15852 14890 15864
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 17696 15892 17724 16136
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16096 18199 16099
rect 18230 16096 18236 16108
rect 18187 16068 18236 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18371 16068 18552 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18524 16040 18552 16068
rect 18506 15988 18512 16040
rect 18564 15988 18570 16040
rect 18616 16028 18644 16136
rect 18708 16096 18736 16204
rect 18782 16192 18788 16244
rect 18840 16192 18846 16244
rect 20901 16235 20959 16241
rect 20901 16201 20913 16235
rect 20947 16201 20959 16235
rect 20901 16195 20959 16201
rect 18800 16164 18828 16192
rect 18800 16136 20760 16164
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 18708 16068 18797 16096
rect 18785 16065 18797 16068
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 19150 16056 19156 16108
rect 19208 16096 19214 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19208 16068 19257 16096
rect 19208 16056 19214 16068
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19521 16099 19579 16105
rect 19521 16065 19533 16099
rect 19567 16096 19579 16099
rect 19610 16096 19616 16108
rect 19567 16068 19616 16096
rect 19567 16065 19579 16068
rect 19521 16059 19579 16065
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19812 16028 19840 16059
rect 20070 16056 20076 16108
rect 20128 16056 20134 16108
rect 18616 16000 19840 16028
rect 19889 16031 19947 16037
rect 19889 15997 19901 16031
rect 19935 16028 19947 16031
rect 20732 16028 20760 16136
rect 20916 16108 20944 16195
rect 21358 16192 21364 16244
rect 21416 16192 21422 16244
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 23566 16232 23572 16244
rect 23339 16204 23572 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 24673 16235 24731 16241
rect 24673 16201 24685 16235
rect 24719 16232 24731 16235
rect 24854 16232 24860 16244
rect 24719 16204 24860 16232
rect 24719 16201 24731 16204
rect 24673 16195 24731 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 21269 16167 21327 16173
rect 21269 16133 21281 16167
rect 21315 16164 21327 16167
rect 22094 16164 22100 16176
rect 21315 16136 22100 16164
rect 21315 16133 21327 16136
rect 21269 16127 21327 16133
rect 22094 16124 22100 16136
rect 22152 16164 22158 16176
rect 22152 16136 23428 16164
rect 22152 16124 22158 16136
rect 20898 16056 20904 16108
rect 20956 16056 20962 16108
rect 22002 16056 22008 16108
rect 22060 16096 22066 16108
rect 23400 16105 23428 16136
rect 25498 16124 25504 16176
rect 25556 16164 25562 16176
rect 26329 16167 26387 16173
rect 26329 16164 26341 16167
rect 25556 16136 26341 16164
rect 25556 16124 25562 16136
rect 26329 16133 26341 16136
rect 26375 16133 26387 16167
rect 26329 16127 26387 16133
rect 23201 16099 23259 16105
rect 23201 16096 23213 16099
rect 22060 16068 23213 16096
rect 22060 16056 22066 16068
rect 23201 16065 23213 16068
rect 23247 16065 23259 16099
rect 23201 16059 23259 16065
rect 23385 16099 23443 16105
rect 23385 16065 23397 16099
rect 23431 16096 23443 16099
rect 23477 16099 23535 16105
rect 23477 16096 23489 16099
rect 23431 16068 23489 16096
rect 23431 16065 23443 16068
rect 23385 16059 23443 16065
rect 23477 16065 23489 16068
rect 23523 16065 23535 16099
rect 23477 16059 23535 16065
rect 23842 16056 23848 16108
rect 23900 16056 23906 16108
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24394 16096 24400 16108
rect 24351 16068 24400 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 26142 16056 26148 16108
rect 26200 16056 26206 16108
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 21453 16031 21511 16037
rect 21453 16028 21465 16031
rect 19935 16000 20116 16028
rect 20732 16000 21465 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 18690 15920 18696 15972
rect 18748 15960 18754 15972
rect 19610 15960 19616 15972
rect 18748 15932 19616 15960
rect 18748 15920 18754 15932
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 20088 15892 20116 16000
rect 21453 15997 21465 16000
rect 21499 16028 21511 16031
rect 22370 16028 22376 16040
rect 21499 16000 22376 16028
rect 21499 15997 21511 16000
rect 21453 15991 21511 15997
rect 22370 15988 22376 16000
rect 22428 15988 22434 16040
rect 24213 16031 24271 16037
rect 24213 15997 24225 16031
rect 24259 15997 24271 16031
rect 26436 16028 26464 16059
rect 26510 16056 26516 16108
rect 26568 16096 26574 16108
rect 27062 16096 27068 16108
rect 26568 16068 27068 16096
rect 26568 16056 26574 16068
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 27522 16028 27528 16040
rect 26436 16000 27528 16028
rect 24213 15991 24271 15997
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 24228 15960 24256 15991
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 23440 15932 24256 15960
rect 23440 15920 23446 15932
rect 25682 15892 25688 15904
rect 17696 15864 25688 15892
rect 25682 15852 25688 15864
rect 25740 15852 25746 15904
rect 26694 15852 26700 15904
rect 26752 15852 26758 15904
rect 1104 15802 31280 15824
rect 1104 15750 4182 15802
rect 4234 15750 4246 15802
rect 4298 15750 4310 15802
rect 4362 15750 4374 15802
rect 4426 15750 4438 15802
rect 4490 15750 4502 15802
rect 4554 15750 10182 15802
rect 10234 15750 10246 15802
rect 10298 15750 10310 15802
rect 10362 15750 10374 15802
rect 10426 15750 10438 15802
rect 10490 15750 10502 15802
rect 10554 15750 16182 15802
rect 16234 15750 16246 15802
rect 16298 15750 16310 15802
rect 16362 15750 16374 15802
rect 16426 15750 16438 15802
rect 16490 15750 16502 15802
rect 16554 15750 22182 15802
rect 22234 15750 22246 15802
rect 22298 15750 22310 15802
rect 22362 15750 22374 15802
rect 22426 15750 22438 15802
rect 22490 15750 22502 15802
rect 22554 15750 28182 15802
rect 28234 15750 28246 15802
rect 28298 15750 28310 15802
rect 28362 15750 28374 15802
rect 28426 15750 28438 15802
rect 28490 15750 28502 15802
rect 28554 15750 31280 15802
rect 1104 15728 31280 15750
rect 1854 15648 1860 15700
rect 1912 15648 1918 15700
rect 3421 15691 3479 15697
rect 3421 15657 3433 15691
rect 3467 15688 3479 15691
rect 4798 15688 4804 15700
rect 3467 15660 4804 15688
rect 3467 15657 3479 15660
rect 3421 15651 3479 15657
rect 4798 15648 4804 15660
rect 4856 15648 4862 15700
rect 6362 15688 6368 15700
rect 5184 15660 6368 15688
rect 1872 15416 1900 15648
rect 2038 15444 2044 15496
rect 2096 15484 2102 15496
rect 5184 15493 5212 15660
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 7892 15660 8309 15688
rect 7892 15648 7898 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 13170 15688 13176 15700
rect 11020 15660 13176 15688
rect 11020 15648 11026 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 13633 15691 13691 15697
rect 13633 15688 13645 15691
rect 13320 15660 13645 15688
rect 13320 15648 13326 15660
rect 13633 15657 13645 15660
rect 13679 15657 13691 15691
rect 13633 15651 13691 15657
rect 11606 15620 11612 15632
rect 10705 15592 11612 15620
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 5169 15487 5227 15493
rect 2096 15456 2774 15484
rect 2096 15444 2102 15456
rect 2286 15419 2344 15425
rect 2286 15416 2298 15419
rect 1872 15388 2298 15416
rect 2286 15385 2298 15388
rect 2332 15385 2344 15419
rect 2746 15416 2774 15456
rect 5169 15453 5181 15487
rect 5215 15453 5227 15487
rect 5169 15447 5227 15453
rect 5445 15487 5503 15493
rect 5445 15453 5457 15487
rect 5491 15484 5503 15487
rect 6917 15487 6975 15493
rect 6917 15484 6929 15487
rect 5491 15456 6929 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 6917 15453 6929 15456
rect 6963 15484 6975 15487
rect 7944 15484 7972 15512
rect 6963 15456 7972 15484
rect 9217 15487 9275 15493
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 10705 15484 10733 15592
rect 11606 15580 11612 15592
rect 11664 15620 11670 15632
rect 11664 15592 12296 15620
rect 11664 15580 11670 15592
rect 10778 15512 10784 15564
rect 10836 15512 10842 15564
rect 10870 15512 10876 15564
rect 10928 15552 10934 15564
rect 12268 15561 12296 15592
rect 11241 15555 11299 15561
rect 11241 15552 11253 15555
rect 10928 15524 11253 15552
rect 10928 15512 10934 15524
rect 11241 15521 11253 15524
rect 11287 15521 11299 15555
rect 11241 15515 11299 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15521 12311 15555
rect 13648 15552 13676 15651
rect 15102 15648 15108 15700
rect 15160 15688 15166 15700
rect 15160 15660 18092 15688
rect 15160 15648 15166 15660
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 16114 15620 16120 15632
rect 15436 15592 16120 15620
rect 15436 15580 15442 15592
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 17957 15623 18015 15629
rect 17957 15589 17969 15623
rect 18003 15589 18015 15623
rect 18064 15620 18092 15660
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 19150 15688 19156 15700
rect 18380 15660 19156 15688
rect 18380 15648 18386 15660
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19426 15648 19432 15700
rect 19484 15648 19490 15700
rect 22646 15688 22652 15700
rect 21008 15660 22652 15688
rect 21008 15620 21036 15660
rect 18064 15592 21036 15620
rect 17957 15583 18015 15589
rect 14645 15555 14703 15561
rect 14645 15552 14657 15555
rect 13648 15524 14657 15552
rect 12253 15515 12311 15521
rect 14645 15521 14657 15524
rect 14691 15521 14703 15555
rect 17972 15552 18000 15583
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 17972 15524 18521 15552
rect 14645 15515 14703 15521
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 18509 15515 18567 15521
rect 18601 15555 18659 15561
rect 18601 15521 18613 15555
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 9263 15456 10733 15484
rect 10796 15484 10824 15512
rect 11422 15484 11428 15496
rect 10796 15456 11428 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 4798 15416 4804 15428
rect 2746 15388 4804 15416
rect 2286 15379 2344 15385
rect 4798 15376 4804 15388
rect 4856 15416 4862 15428
rect 5460 15416 5488 15447
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 4856 15388 5488 15416
rect 5712 15419 5770 15425
rect 4856 15376 4862 15388
rect 5712 15385 5724 15419
rect 5758 15416 5770 15419
rect 5810 15416 5816 15428
rect 5758 15388 5816 15416
rect 5758 15385 5770 15388
rect 5712 15379 5770 15385
rect 5810 15376 5816 15388
rect 5868 15376 5874 15428
rect 7162 15419 7220 15425
rect 7162 15416 7174 15419
rect 6288 15388 7174 15416
rect 5353 15351 5411 15357
rect 5353 15317 5365 15351
rect 5399 15348 5411 15351
rect 6288 15348 6316 15388
rect 7162 15385 7174 15388
rect 7208 15385 7220 15419
rect 7162 15379 7220 15385
rect 9484 15419 9542 15425
rect 9484 15385 9496 15419
rect 9530 15416 9542 15419
rect 9582 15416 9588 15428
rect 9530 15388 9588 15416
rect 9530 15385 9542 15388
rect 9484 15379 9542 15385
rect 9582 15376 9588 15388
rect 9640 15376 9646 15428
rect 11882 15416 11888 15428
rect 10612 15388 11888 15416
rect 5399 15320 6316 15348
rect 6825 15351 6883 15357
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 6825 15317 6837 15351
rect 6871 15348 6883 15351
rect 7742 15348 7748 15360
rect 6871 15320 7748 15348
rect 6871 15317 6883 15320
rect 6825 15311 6883 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 10612 15357 10640 15388
rect 11882 15376 11888 15388
rect 11940 15416 11946 15428
rect 12084 15416 12112 15447
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12509 15487 12567 15493
rect 12509 15484 12521 15487
rect 12216 15456 12521 15484
rect 12216 15444 12222 15456
rect 12509 15453 12521 15456
rect 12555 15453 12567 15487
rect 12509 15447 12567 15453
rect 15562 15444 15568 15496
rect 15620 15484 15626 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15620 15456 15853 15484
rect 15620 15444 15626 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 15841 15447 15899 15453
rect 16224 15456 17693 15484
rect 11940 15388 12112 15416
rect 11940 15376 11946 15388
rect 16224 15360 16252 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 17773 15487 17831 15493
rect 17773 15453 17785 15487
rect 17819 15484 17831 15487
rect 18322 15484 18328 15496
rect 17819 15456 18328 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 17696 15416 17724 15447
rect 18322 15444 18328 15456
rect 18380 15444 18386 15496
rect 18616 15484 18644 15515
rect 20898 15512 20904 15564
rect 20956 15512 20962 15564
rect 22572 15552 22600 15660
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 23017 15691 23075 15697
rect 23017 15657 23029 15691
rect 23063 15688 23075 15691
rect 23842 15688 23848 15700
rect 23063 15660 23848 15688
rect 23063 15657 23075 15660
rect 23017 15651 23075 15657
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 26694 15648 26700 15700
rect 26752 15648 26758 15700
rect 27522 15648 27528 15700
rect 27580 15688 27586 15700
rect 28537 15691 28595 15697
rect 28537 15688 28549 15691
rect 27580 15660 28549 15688
rect 27580 15648 27586 15660
rect 28537 15657 28549 15660
rect 28583 15657 28595 15691
rect 28537 15651 28595 15657
rect 25866 15552 25872 15564
rect 22572 15524 25872 15552
rect 25866 15512 25872 15524
rect 25924 15512 25930 15564
rect 26712 15552 26740 15648
rect 28353 15555 28411 15561
rect 28353 15552 28365 15555
rect 26712 15524 28365 15552
rect 28353 15521 28365 15524
rect 28399 15521 28411 15555
rect 28353 15515 28411 15521
rect 29181 15555 29239 15561
rect 29181 15521 29193 15555
rect 29227 15552 29239 15555
rect 29638 15552 29644 15564
rect 29227 15524 29644 15552
rect 29227 15521 29239 15524
rect 29181 15515 29239 15521
rect 29638 15512 29644 15524
rect 29696 15512 29702 15564
rect 19702 15484 19708 15496
rect 18524 15456 18644 15484
rect 19516 15459 19708 15484
rect 19475 15456 19708 15459
rect 18524 15428 18552 15456
rect 19475 15453 19544 15456
rect 17862 15416 17868 15428
rect 17696 15388 17868 15416
rect 17862 15376 17868 15388
rect 17920 15376 17926 15428
rect 17957 15419 18015 15425
rect 17957 15385 17969 15419
rect 18003 15416 18015 15419
rect 18003 15388 18460 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 10597 15351 10655 15357
rect 10597 15317 10609 15351
rect 10643 15317 10655 15351
rect 10597 15311 10655 15317
rect 10686 15308 10692 15360
rect 10744 15308 10750 15360
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 11020 15320 11069 15348
rect 11020 15308 11026 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 11149 15351 11207 15357
rect 11149 15317 11161 15351
rect 11195 15348 11207 15351
rect 11517 15351 11575 15357
rect 11517 15348 11529 15351
rect 11195 15320 11529 15348
rect 11195 15317 11207 15320
rect 11149 15311 11207 15317
rect 11517 15317 11529 15320
rect 11563 15317 11575 15351
rect 11517 15311 11575 15317
rect 14090 15308 14096 15360
rect 14148 15308 14154 15360
rect 15286 15308 15292 15360
rect 15344 15308 15350 15360
rect 16206 15308 16212 15360
rect 16264 15308 16270 15360
rect 18046 15308 18052 15360
rect 18104 15308 18110 15360
rect 18432 15357 18460 15388
rect 18506 15376 18512 15428
rect 18564 15376 18570 15428
rect 19242 15376 19248 15428
rect 19300 15376 19306 15428
rect 19475 15419 19487 15453
rect 19521 15422 19544 15453
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 20916 15484 20944 15512
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 20916 15456 21005 15484
rect 20993 15453 21005 15456
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 26050 15444 26056 15496
rect 26108 15444 26114 15496
rect 26510 15444 26516 15496
rect 26568 15484 26574 15496
rect 27709 15487 27767 15493
rect 27709 15484 27721 15487
rect 26568 15456 27721 15484
rect 26568 15444 26574 15456
rect 27709 15453 27721 15456
rect 27755 15453 27767 15487
rect 27709 15447 27767 15453
rect 19521 15419 19533 15422
rect 19475 15413 19533 15419
rect 21545 15419 21603 15425
rect 21545 15416 21557 15419
rect 21192 15388 21557 15416
rect 18417 15351 18475 15357
rect 18417 15317 18429 15351
rect 18463 15348 18475 15351
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 18463 15320 19625 15348
rect 18463 15317 18475 15320
rect 18417 15311 18475 15317
rect 19613 15317 19625 15320
rect 19659 15348 19671 15351
rect 20530 15348 20536 15360
rect 19659 15320 20536 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 21192 15357 21220 15388
rect 21545 15385 21557 15388
rect 21591 15385 21603 15419
rect 21545 15379 21603 15385
rect 22002 15376 22008 15428
rect 22060 15376 22066 15428
rect 24118 15376 24124 15428
rect 24176 15416 24182 15428
rect 26881 15419 26939 15425
rect 26881 15416 26893 15419
rect 24176 15388 26893 15416
rect 24176 15376 24182 15388
rect 26881 15385 26893 15388
rect 26927 15416 26939 15419
rect 26970 15416 26976 15428
rect 26927 15388 26976 15416
rect 26927 15385 26939 15388
rect 26881 15379 26939 15385
rect 26970 15376 26976 15388
rect 27028 15416 27034 15428
rect 27430 15416 27436 15428
rect 27028 15388 27436 15416
rect 27028 15376 27034 15388
rect 27430 15376 27436 15388
rect 27488 15376 27494 15428
rect 21177 15351 21235 15357
rect 21177 15317 21189 15351
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 26694 15308 26700 15360
rect 26752 15308 26758 15360
rect 27798 15308 27804 15360
rect 27856 15308 27862 15360
rect 1104 15258 31280 15280
rect 1104 15206 4922 15258
rect 4974 15206 4986 15258
rect 5038 15206 5050 15258
rect 5102 15206 5114 15258
rect 5166 15206 5178 15258
rect 5230 15206 5242 15258
rect 5294 15206 10922 15258
rect 10974 15206 10986 15258
rect 11038 15206 11050 15258
rect 11102 15206 11114 15258
rect 11166 15206 11178 15258
rect 11230 15206 11242 15258
rect 11294 15206 16922 15258
rect 16974 15206 16986 15258
rect 17038 15206 17050 15258
rect 17102 15206 17114 15258
rect 17166 15206 17178 15258
rect 17230 15206 17242 15258
rect 17294 15206 22922 15258
rect 22974 15206 22986 15258
rect 23038 15206 23050 15258
rect 23102 15206 23114 15258
rect 23166 15206 23178 15258
rect 23230 15206 23242 15258
rect 23294 15206 28922 15258
rect 28974 15206 28986 15258
rect 29038 15206 29050 15258
rect 29102 15206 29114 15258
rect 29166 15206 29178 15258
rect 29230 15206 29242 15258
rect 29294 15206 31280 15258
rect 1104 15184 31280 15206
rect 5810 15104 5816 15156
rect 5868 15104 5874 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 6825 15147 6883 15153
rect 6825 15144 6837 15147
rect 6696 15116 6837 15144
rect 6696 15104 6702 15116
rect 6825 15113 6837 15116
rect 6871 15113 6883 15147
rect 6825 15107 6883 15113
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 7892 15116 8156 15144
rect 7892 15104 7898 15116
rect 7300 15048 7972 15076
rect 7300 15020 7328 15048
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 15008 6055 15011
rect 6733 15011 6791 15017
rect 6043 14980 6408 15008
rect 6043 14977 6055 14980
rect 5997 14971 6055 14977
rect 6380 14881 6408 14980
rect 6733 14977 6745 15011
rect 6779 15008 6791 15011
rect 7193 15011 7251 15017
rect 7193 15008 7205 15011
rect 6779 14980 7205 15008
rect 6779 14977 6791 14980
rect 6733 14971 6791 14977
rect 7193 14977 7205 14980
rect 7239 14977 7251 15011
rect 7193 14971 7251 14977
rect 7282 14968 7288 15020
rect 7340 14968 7346 15020
rect 7742 14968 7748 15020
rect 7800 14968 7806 15020
rect 7944 15017 7972 15048
rect 8128 15017 8156 15116
rect 9582 15104 9588 15156
rect 9640 15104 9646 15156
rect 10686 15104 10692 15156
rect 10744 15104 10750 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13170 15104 13176 15156
rect 13228 15104 13234 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 14090 15144 14096 15156
rect 13311 15116 14096 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14458 15104 14464 15156
rect 14516 15144 14522 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 14516 15116 14933 15144
rect 14516 15104 14522 15116
rect 14921 15113 14933 15116
rect 14967 15113 14979 15147
rect 14921 15107 14979 15113
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15286 15144 15292 15156
rect 15059 15116 15292 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 15930 15104 15936 15156
rect 15988 15144 15994 15156
rect 16485 15147 16543 15153
rect 16485 15144 16497 15147
rect 15988 15116 16497 15144
rect 15988 15104 15994 15116
rect 16485 15113 16497 15116
rect 16531 15113 16543 15147
rect 16485 15107 16543 15113
rect 18046 15104 18052 15156
rect 18104 15104 18110 15156
rect 21913 15147 21971 15153
rect 21913 15113 21925 15147
rect 21959 15144 21971 15147
rect 22002 15144 22008 15156
rect 21959 15116 22008 15144
rect 21959 15113 21971 15116
rect 21913 15107 21971 15113
rect 22002 15104 22008 15116
rect 22060 15104 22066 15156
rect 25501 15147 25559 15153
rect 25501 15113 25513 15147
rect 25547 15144 25559 15147
rect 26142 15144 26148 15156
rect 25547 15116 26148 15144
rect 25547 15113 25559 15116
rect 25501 15107 25559 15113
rect 26142 15104 26148 15116
rect 26200 15104 26206 15156
rect 26329 15147 26387 15153
rect 26329 15113 26341 15147
rect 26375 15144 26387 15147
rect 26694 15144 26700 15156
rect 26375 15116 26700 15144
rect 26375 15113 26387 15116
rect 26329 15107 26387 15113
rect 26694 15104 26700 15116
rect 26752 15104 26758 15156
rect 26789 15147 26847 15153
rect 26789 15113 26801 15147
rect 26835 15113 26847 15147
rect 26789 15107 26847 15113
rect 8202 15036 8208 15088
rect 8260 15036 8266 15088
rect 8478 15017 8484 15020
rect 7929 15011 7987 15017
rect 7929 14977 7941 15011
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 8077 15011 8156 15017
rect 8077 14977 8089 15011
rect 8123 14980 8156 15011
rect 8297 15011 8355 15017
rect 8123 14977 8135 14980
rect 8077 14971 8135 14977
rect 8297 14977 8309 15011
rect 8343 14977 8355 15011
rect 8297 14971 8355 14977
rect 8435 15011 8484 15017
rect 8435 14977 8447 15011
rect 8481 14977 8484 15011
rect 8435 14971 8484 14977
rect 6917 14943 6975 14949
rect 6917 14940 6929 14943
rect 6748 14912 6929 14940
rect 6748 14884 6776 14912
rect 6917 14909 6929 14912
rect 6963 14909 6975 14943
rect 7760 14940 7788 14968
rect 8312 14940 8340 14971
rect 8478 14968 8484 14971
rect 8536 14968 8542 15020
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 10704 15008 10732 15104
rect 16206 15076 16212 15088
rect 11716 15048 16212 15076
rect 11716 15020 11744 15048
rect 9815 14980 10732 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 12636 14980 14688 15008
rect 7760 14912 8340 14940
rect 6917 14903 6975 14909
rect 12434 14900 12440 14952
rect 12492 14900 12498 14952
rect 6365 14875 6423 14881
rect 6365 14841 6377 14875
rect 6411 14841 6423 14875
rect 6365 14835 6423 14841
rect 6730 14832 6736 14884
rect 6788 14832 6794 14884
rect 7282 14832 7288 14884
rect 7340 14872 7346 14884
rect 8202 14872 8208 14884
rect 7340 14844 8208 14872
rect 7340 14832 7346 14844
rect 8202 14832 8208 14844
rect 8260 14832 8266 14884
rect 8573 14875 8631 14881
rect 8573 14841 8585 14875
rect 8619 14872 8631 14875
rect 12636 14872 12664 14980
rect 13446 14900 13452 14952
rect 13504 14900 13510 14952
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13688 14912 14197 14940
rect 13688 14900 13694 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 8619 14844 12664 14872
rect 12728 14844 13676 14872
rect 8619 14841 8631 14844
rect 8573 14835 8631 14841
rect 11882 14764 11888 14816
rect 11940 14764 11946 14816
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12728 14804 12756 14844
rect 13648 14813 13676 14844
rect 12216 14776 12756 14804
rect 13633 14807 13691 14813
rect 12216 14764 12222 14776
rect 13633 14773 13645 14807
rect 13679 14773 13691 14807
rect 13633 14767 13691 14773
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 13780 14776 14565 14804
rect 13780 14764 13786 14776
rect 14553 14773 14565 14776
rect 14599 14773 14611 14807
rect 14660 14804 14688 14980
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15562 15017 15568 15020
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15252 14980 15393 15008
rect 15252 14968 15258 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 15529 15011 15568 15017
rect 15529 14977 15541 15011
rect 15529 14971 15568 14977
rect 15562 14968 15568 14971
rect 15620 14968 15626 15020
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 15746 14968 15752 15020
rect 15804 14968 15810 15020
rect 15861 15017 15889 15048
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 15846 15011 15904 15017
rect 15846 14977 15858 15011
rect 15892 14977 15904 15011
rect 15846 14971 15904 14977
rect 16114 14968 16120 15020
rect 16172 14968 16178 15020
rect 17681 15011 17739 15017
rect 17681 14977 17693 15011
rect 17727 15008 17739 15011
rect 18064 15008 18092 15104
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 17727 14980 18092 15008
rect 18156 14980 18613 15008
rect 17727 14977 17739 14980
rect 17681 14971 17739 14977
rect 14734 14900 14740 14952
rect 14792 14940 14798 14952
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 14792 14912 15117 14940
rect 14792 14900 14798 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 15672 14940 15700 14968
rect 16209 14943 16267 14949
rect 16209 14940 16221 14943
rect 15105 14903 15163 14909
rect 15304 14912 15700 14940
rect 16040 14912 16221 14940
rect 15304 14884 15332 14912
rect 15286 14832 15292 14884
rect 15344 14832 15350 14884
rect 16040 14881 16068 14912
rect 16209 14909 16221 14912
rect 16255 14909 16267 14943
rect 16209 14903 16267 14909
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 18156 14940 18184 14980
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 18785 15011 18843 15017
rect 18785 14977 18797 15011
rect 18831 15008 18843 15011
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18831 14980 18889 15008
rect 18831 14977 18843 14980
rect 18785 14971 18843 14977
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 17920 14912 18184 14940
rect 18417 14943 18475 14949
rect 17920 14900 17926 14912
rect 18417 14909 18429 14943
rect 18463 14940 18475 14943
rect 18506 14940 18512 14952
rect 18463 14912 18512 14940
rect 18463 14909 18475 14912
rect 18417 14903 18475 14909
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 18616 14940 18644 14971
rect 20530 14968 20536 15020
rect 20588 14968 20594 15020
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 21910 15008 21916 15020
rect 21315 14980 21916 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22002 14968 22008 15020
rect 22060 14968 22066 15020
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 23842 15008 23848 15020
rect 22888 14980 23848 15008
rect 22888 14968 22894 14980
rect 23842 14968 23848 14980
rect 23900 14968 23906 15020
rect 25682 14968 25688 15020
rect 25740 15008 25746 15020
rect 26142 15008 26148 15020
rect 25740 14980 26148 15008
rect 25740 14968 25746 14980
rect 26142 14968 26148 14980
rect 26200 14968 26206 15020
rect 26418 14968 26424 15020
rect 26476 15008 26482 15020
rect 26804 15008 26832 15107
rect 27246 15104 27252 15156
rect 27304 15104 27310 15156
rect 29181 15147 29239 15153
rect 29181 15113 29193 15147
rect 29227 15144 29239 15147
rect 29638 15144 29644 15156
rect 29227 15116 29644 15144
rect 29227 15113 29239 15116
rect 29181 15107 29239 15113
rect 29638 15104 29644 15116
rect 29696 15104 29702 15156
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26476 14980 26556 15008
rect 26804 14980 26985 15008
rect 26476 14968 26482 14980
rect 24302 14940 24308 14952
rect 18616 14912 24308 14940
rect 24302 14900 24308 14912
rect 24360 14900 24366 14952
rect 25961 14943 26019 14949
rect 25961 14909 25973 14943
rect 26007 14940 26019 14943
rect 26050 14940 26056 14952
rect 26007 14912 26056 14940
rect 26007 14909 26019 14912
rect 25961 14903 26019 14909
rect 26050 14900 26056 14912
rect 26108 14900 26114 14952
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14940 26295 14943
rect 26326 14940 26332 14952
rect 26283 14912 26332 14940
rect 26283 14909 26295 14912
rect 26237 14903 26295 14909
rect 26326 14900 26332 14912
rect 26384 14900 26390 14952
rect 26528 14940 26556 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 27264 15008 27292 15104
rect 27709 15079 27767 15085
rect 27709 15045 27721 15079
rect 27755 15076 27767 15079
rect 27798 15076 27804 15088
rect 27755 15048 27804 15076
rect 27755 15045 27767 15048
rect 27709 15039 27767 15045
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 29365 15079 29423 15085
rect 29365 15076 29377 15079
rect 28934 15048 29377 15076
rect 29365 15045 29377 15048
rect 29411 15045 29423 15079
rect 29365 15039 29423 15045
rect 26973 14971 27031 14977
rect 27080 14980 27292 15008
rect 29457 15011 29515 15017
rect 27080 14940 27108 14980
rect 29457 14977 29469 15011
rect 29503 14977 29515 15011
rect 29457 14971 29515 14977
rect 26528 14912 27108 14940
rect 27154 14900 27160 14952
rect 27212 14940 27218 14952
rect 27433 14943 27491 14949
rect 27433 14940 27445 14943
rect 27212 14912 27445 14940
rect 27212 14900 27218 14912
rect 27433 14909 27445 14912
rect 27479 14909 27491 14943
rect 29362 14940 29368 14952
rect 27433 14903 27491 14909
rect 27540 14912 29368 14940
rect 16025 14875 16083 14881
rect 16025 14841 16037 14875
rect 16071 14841 16083 14875
rect 16025 14835 16083 14841
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 22002 14872 22008 14884
rect 18012 14844 22008 14872
rect 18012 14832 18018 14844
rect 22002 14832 22008 14844
rect 22060 14872 22066 14884
rect 26510 14872 26516 14884
rect 22060 14844 26516 14872
rect 22060 14832 22066 14844
rect 26510 14832 26516 14844
rect 26568 14872 26574 14884
rect 27540 14872 27568 14912
rect 29362 14900 29368 14912
rect 29420 14940 29426 14952
rect 29472 14940 29500 14971
rect 29420 14912 29500 14940
rect 29420 14900 29426 14912
rect 26568 14844 27568 14872
rect 26568 14832 26574 14844
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 14660 14776 16129 14804
rect 14553 14767 14611 14773
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 16117 14767 16175 14773
rect 17494 14764 17500 14816
rect 17552 14764 17558 14816
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 19024 14776 19073 14804
rect 19024 14764 19030 14776
rect 19061 14773 19073 14776
rect 19107 14804 19119 14807
rect 19334 14804 19340 14816
rect 19107 14776 19340 14804
rect 19107 14773 19119 14776
rect 19061 14767 19119 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 24670 14804 24676 14816
rect 20680 14776 24676 14804
rect 20680 14764 20686 14776
rect 24670 14764 24676 14776
rect 24728 14764 24734 14816
rect 25866 14764 25872 14816
rect 25924 14804 25930 14816
rect 26786 14804 26792 14816
rect 25924 14776 26792 14804
rect 25924 14764 25930 14776
rect 26786 14764 26792 14776
rect 26844 14764 26850 14816
rect 27157 14807 27215 14813
rect 27157 14773 27169 14807
rect 27203 14804 27215 14807
rect 27246 14804 27252 14816
rect 27203 14776 27252 14804
rect 27203 14773 27215 14776
rect 27157 14767 27215 14773
rect 27246 14764 27252 14776
rect 27304 14764 27310 14816
rect 1104 14714 31280 14736
rect 1104 14662 4182 14714
rect 4234 14662 4246 14714
rect 4298 14662 4310 14714
rect 4362 14662 4374 14714
rect 4426 14662 4438 14714
rect 4490 14662 4502 14714
rect 4554 14662 10182 14714
rect 10234 14662 10246 14714
rect 10298 14662 10310 14714
rect 10362 14662 10374 14714
rect 10426 14662 10438 14714
rect 10490 14662 10502 14714
rect 10554 14662 16182 14714
rect 16234 14662 16246 14714
rect 16298 14662 16310 14714
rect 16362 14662 16374 14714
rect 16426 14662 16438 14714
rect 16490 14662 16502 14714
rect 16554 14662 22182 14714
rect 22234 14662 22246 14714
rect 22298 14662 22310 14714
rect 22362 14662 22374 14714
rect 22426 14662 22438 14714
rect 22490 14662 22502 14714
rect 22554 14662 28182 14714
rect 28234 14662 28246 14714
rect 28298 14662 28310 14714
rect 28362 14662 28374 14714
rect 28426 14662 28438 14714
rect 28490 14662 28502 14714
rect 28554 14662 31280 14714
rect 1104 14640 31280 14662
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 15286 14600 15292 14612
rect 11480 14572 15292 14600
rect 11480 14560 11486 14572
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 15562 14560 15568 14612
rect 15620 14560 15626 14612
rect 17586 14600 17592 14612
rect 15672 14572 17592 14600
rect 13906 14492 13912 14544
rect 13964 14492 13970 14544
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 11882 14424 11888 14476
rect 11940 14424 11946 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13504 14436 14320 14464
rect 13504 14424 13510 14436
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 13541 14331 13599 14337
rect 13541 14328 13553 14331
rect 13110 14300 13553 14328
rect 13541 14297 13553 14300
rect 13587 14297 13599 14331
rect 13648 14328 13676 14359
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 14182 14356 14188 14408
rect 14240 14356 14246 14408
rect 14292 14396 14320 14436
rect 15672 14396 15700 14572
rect 17586 14560 17592 14572
rect 17644 14600 17650 14612
rect 17644 14572 18184 14600
rect 17644 14560 17650 14572
rect 18156 14532 18184 14572
rect 18506 14560 18512 14612
rect 18564 14600 18570 14612
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 18564 14572 18613 14600
rect 18564 14560 18570 14572
rect 18601 14569 18613 14572
rect 18647 14569 18659 14603
rect 18601 14563 18659 14569
rect 26050 14560 26056 14612
rect 26108 14600 26114 14612
rect 26329 14603 26387 14609
rect 26329 14600 26341 14603
rect 26108 14572 26341 14600
rect 26108 14560 26114 14572
rect 26329 14569 26341 14572
rect 26375 14569 26387 14603
rect 26329 14563 26387 14569
rect 18156 14504 22094 14532
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17494 14464 17500 14476
rect 17175 14436 17500 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 22066 14464 22094 14504
rect 26326 14464 26332 14476
rect 22066 14436 26332 14464
rect 26326 14424 26332 14436
rect 26384 14424 26390 14476
rect 14292 14368 15700 14396
rect 16850 14356 16856 14408
rect 16908 14356 16914 14408
rect 26234 14356 26240 14408
rect 26292 14396 26298 14408
rect 27154 14396 27160 14408
rect 26292 14368 27160 14396
rect 26292 14356 26298 14368
rect 27154 14356 27160 14368
rect 27212 14396 27218 14408
rect 27709 14399 27767 14405
rect 27709 14396 27721 14399
rect 27212 14368 27721 14396
rect 27212 14356 27218 14368
rect 27709 14365 27721 14368
rect 27755 14365 27767 14399
rect 27709 14359 27767 14365
rect 13648 14300 13768 14328
rect 13541 14291 13599 14297
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13357 14263 13415 14269
rect 13357 14260 13369 14263
rect 13320 14232 13369 14260
rect 13320 14220 13326 14232
rect 13357 14229 13369 14232
rect 13403 14260 13415 14263
rect 13630 14260 13636 14272
rect 13403 14232 13636 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 13740 14260 13768 14300
rect 13906 14288 13912 14340
rect 13964 14328 13970 14340
rect 14430 14331 14488 14337
rect 14430 14328 14442 14331
rect 13964 14300 14442 14328
rect 13964 14288 13970 14300
rect 14430 14297 14442 14300
rect 14476 14297 14488 14331
rect 14430 14291 14488 14297
rect 17862 14288 17868 14340
rect 17920 14288 17926 14340
rect 27246 14288 27252 14340
rect 27304 14328 27310 14340
rect 27442 14331 27500 14337
rect 27442 14328 27454 14331
rect 27304 14300 27454 14328
rect 27304 14288 27310 14300
rect 27442 14297 27454 14300
rect 27488 14297 27500 14331
rect 27442 14291 27500 14297
rect 17954 14260 17960 14272
rect 13740 14232 17960 14260
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 1104 14170 31280 14192
rect 1104 14118 4922 14170
rect 4974 14118 4986 14170
rect 5038 14118 5050 14170
rect 5102 14118 5114 14170
rect 5166 14118 5178 14170
rect 5230 14118 5242 14170
rect 5294 14118 10922 14170
rect 10974 14118 10986 14170
rect 11038 14118 11050 14170
rect 11102 14118 11114 14170
rect 11166 14118 11178 14170
rect 11230 14118 11242 14170
rect 11294 14118 16922 14170
rect 16974 14118 16986 14170
rect 17038 14118 17050 14170
rect 17102 14118 17114 14170
rect 17166 14118 17178 14170
rect 17230 14118 17242 14170
rect 17294 14118 22922 14170
rect 22974 14118 22986 14170
rect 23038 14118 23050 14170
rect 23102 14118 23114 14170
rect 23166 14118 23178 14170
rect 23230 14118 23242 14170
rect 23294 14118 28922 14170
rect 28974 14118 28986 14170
rect 29038 14118 29050 14170
rect 29102 14118 29114 14170
rect 29166 14118 29178 14170
rect 29230 14118 29242 14170
rect 29294 14118 31280 14170
rect 1104 14096 31280 14118
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 4062 14056 4068 14068
rect 3108 14028 4068 14056
rect 3108 14016 3114 14028
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 8849 14059 8907 14065
rect 8849 14025 8861 14059
rect 8895 14056 8907 14059
rect 8938 14056 8944 14068
rect 8895 14028 8944 14056
rect 8895 14025 8907 14028
rect 8849 14019 8907 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 12434 14056 12440 14068
rect 11931 14028 12440 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 12158 13948 12164 14000
rect 12216 13948 12222 14000
rect 12250 13948 12256 14000
rect 12308 13948 12314 14000
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 14292 13988 14320 14019
rect 15746 14016 15752 14068
rect 15804 14016 15810 14068
rect 17862 14016 17868 14068
rect 17920 14016 17926 14068
rect 24765 14059 24823 14065
rect 24765 14025 24777 14059
rect 24811 14056 24823 14059
rect 25498 14056 25504 14068
rect 24811 14028 25504 14056
rect 24811 14025 24823 14028
rect 24765 14019 24823 14025
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 14614 13991 14672 13997
rect 14614 13988 14626 13991
rect 12400 13960 14228 13988
rect 14292 13960 14626 13988
rect 12400 13948 12406 13960
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2866 13920 2872 13932
rect 2547 13892 2872 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 2961 13923 3019 13929
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 3007 13892 3433 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 3421 13889 3433 13892
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 12069 13923 12127 13929
rect 12069 13889 12081 13923
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 3145 13855 3203 13861
rect 3145 13821 3157 13855
rect 3191 13852 3203 13855
rect 3234 13852 3240 13864
rect 3191 13824 3240 13852
rect 3191 13821 3203 13824
rect 3145 13815 3203 13821
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 8478 13784 8484 13796
rect 7892 13756 8484 13784
rect 7892 13744 7898 13756
rect 8478 13744 8484 13756
rect 8536 13744 8542 13796
rect 8680 13728 8708 13883
rect 9674 13812 9680 13864
rect 9732 13812 9738 13864
rect 12084 13852 12112 13883
rect 12360 13852 12388 13948
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12802 13920 12808 13932
rect 12483 13892 12808 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14200 13920 14228 13960
rect 14614 13957 14626 13960
rect 14660 13957 14672 13991
rect 18690 13988 18696 14000
rect 14614 13951 14672 13957
rect 15028 13960 18696 13988
rect 15028 13920 15056 13960
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 14200 13892 15056 13920
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15160 13892 15700 13920
rect 15160 13880 15166 13892
rect 12084 13824 12388 13852
rect 14182 13812 14188 13864
rect 14240 13852 14246 13864
rect 14369 13855 14427 13861
rect 14369 13852 14381 13855
rect 14240 13824 14381 13852
rect 14240 13812 14246 13824
rect 14369 13821 14381 13824
rect 14415 13821 14427 13855
rect 15672 13852 15700 13892
rect 15746 13880 15752 13932
rect 15804 13920 15810 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 15804 13892 16405 13920
rect 15804 13880 15810 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 17773 13923 17831 13929
rect 17773 13889 17785 13923
rect 17819 13920 17831 13923
rect 24118 13920 24124 13932
rect 17819 13892 24124 13920
rect 17819 13889 17831 13892
rect 17773 13883 17831 13889
rect 17788 13852 17816 13883
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24394 13880 24400 13932
rect 24452 13880 24458 13932
rect 15672 13824 17816 13852
rect 14369 13815 14427 13821
rect 24210 13812 24216 13864
rect 24268 13852 24274 13864
rect 24489 13855 24547 13861
rect 24489 13852 24501 13855
rect 24268 13824 24501 13852
rect 24268 13812 24274 13824
rect 24489 13821 24501 13824
rect 24535 13821 24547 13855
rect 24489 13815 24547 13821
rect 2222 13676 2228 13728
rect 2280 13716 2286 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 2280 13688 2329 13716
rect 2280 13676 2286 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2317 13679 2375 13685
rect 2590 13676 2596 13728
rect 2648 13676 2654 13728
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 8662 13716 8668 13728
rect 4212 13688 8668 13716
rect 4212 13676 4218 13688
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9122 13676 9128 13728
rect 9180 13676 9186 13728
rect 15838 13676 15844 13728
rect 15896 13676 15902 13728
rect 21358 13676 21364 13728
rect 21416 13716 21422 13728
rect 24397 13719 24455 13725
rect 24397 13716 24409 13719
rect 21416 13688 24409 13716
rect 21416 13676 21422 13688
rect 24397 13685 24409 13688
rect 24443 13685 24455 13719
rect 24397 13679 24455 13685
rect 1104 13626 31280 13648
rect 1104 13574 4182 13626
rect 4234 13574 4246 13626
rect 4298 13574 4310 13626
rect 4362 13574 4374 13626
rect 4426 13574 4438 13626
rect 4490 13574 4502 13626
rect 4554 13574 10182 13626
rect 10234 13574 10246 13626
rect 10298 13574 10310 13626
rect 10362 13574 10374 13626
rect 10426 13574 10438 13626
rect 10490 13574 10502 13626
rect 10554 13574 16182 13626
rect 16234 13574 16246 13626
rect 16298 13574 16310 13626
rect 16362 13574 16374 13626
rect 16426 13574 16438 13626
rect 16490 13574 16502 13626
rect 16554 13574 22182 13626
rect 22234 13574 22246 13626
rect 22298 13574 22310 13626
rect 22362 13574 22374 13626
rect 22426 13574 22438 13626
rect 22490 13574 22502 13626
rect 22554 13574 28182 13626
rect 28234 13574 28246 13626
rect 28298 13574 28310 13626
rect 28362 13574 28374 13626
rect 28426 13574 28438 13626
rect 28490 13574 28502 13626
rect 28554 13574 31280 13626
rect 1104 13552 31280 13574
rect 2590 13512 2596 13524
rect 1688 13484 2596 13512
rect 1688 13317 1716 13484
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 2924 13484 3801 13512
rect 2924 13472 2930 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 4154 13472 4160 13524
rect 4212 13472 4218 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4706 13512 4712 13524
rect 4580 13484 4712 13512
rect 4580 13472 4586 13484
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 7742 13512 7748 13524
rect 7116 13484 7748 13512
rect 3329 13447 3387 13453
rect 3329 13413 3341 13447
rect 3375 13444 3387 13447
rect 3988 13444 4016 13472
rect 3375 13416 4016 13444
rect 3375 13413 3387 13416
rect 3329 13407 3387 13413
rect 4172 13376 4200 13472
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4172 13348 4261 13376
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4614 13376 4620 13388
rect 4479 13348 4620 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6012 13348 6561 13376
rect 6012 13320 6040 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2038 13308 2044 13320
rect 1995 13280 2044 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2038 13268 2044 13280
rect 2096 13268 2102 13320
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 3844 13280 5181 13308
rect 3844 13268 3850 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5994 13317 6000 13320
rect 5813 13311 5871 13317
rect 5813 13277 5825 13311
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5961 13311 6000 13317
rect 5961 13277 5973 13311
rect 5961 13271 6000 13277
rect 2194 13243 2252 13249
rect 2194 13240 2206 13243
rect 1872 13212 2206 13240
rect 1872 13181 1900 13212
rect 2194 13209 2206 13212
rect 2240 13209 2252 13243
rect 2194 13203 2252 13209
rect 4157 13243 4215 13249
rect 4157 13209 4169 13243
rect 4203 13240 4215 13243
rect 4617 13243 4675 13249
rect 4617 13240 4629 13243
rect 4203 13212 4629 13240
rect 4203 13209 4215 13212
rect 4157 13203 4215 13209
rect 4617 13209 4629 13212
rect 4663 13209 4675 13243
rect 4617 13203 4675 13209
rect 4706 13200 4712 13252
rect 4764 13240 4770 13252
rect 5828 13240 5856 13271
rect 5994 13268 6000 13271
rect 6052 13268 6058 13320
rect 6319 13311 6377 13317
rect 6319 13277 6331 13311
rect 6365 13308 6377 13311
rect 7116 13308 7144 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9674 13512 9680 13524
rect 8803 13484 9680 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14148 13484 14841 13512
rect 14148 13472 14154 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 14829 13475 14887 13481
rect 15470 13472 15476 13524
rect 15528 13512 15534 13524
rect 16114 13512 16120 13524
rect 15528 13484 16120 13512
rect 15528 13472 15534 13484
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 25866 13512 25872 13524
rect 22572 13484 25872 13512
rect 9582 13404 9588 13456
rect 9640 13404 9646 13456
rect 9692 13444 9720 13472
rect 20622 13444 20628 13456
rect 9692 13416 10088 13444
rect 8662 13336 8668 13388
rect 8720 13376 8726 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 8720 13348 9413 13376
rect 8720 13336 8726 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 9600 13376 9628 13404
rect 9950 13376 9956 13388
rect 9539 13348 9956 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 6365 13280 7144 13308
rect 6365 13277 6377 13280
rect 6319 13271 6377 13277
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7374 13268 7380 13320
rect 7432 13268 7438 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 9309 13311 9367 13317
rect 9309 13308 9321 13311
rect 9180 13280 9321 13308
rect 9180 13268 9186 13280
rect 9309 13277 9321 13280
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 4764 13212 5856 13240
rect 6089 13243 6147 13249
rect 4764 13200 4770 13212
rect 6089 13209 6101 13243
rect 6135 13209 6147 13243
rect 6089 13203 6147 13209
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 5350 13132 5356 13184
rect 5408 13132 5414 13184
rect 6104 13172 6132 13203
rect 6178 13200 6184 13252
rect 6236 13200 6242 13252
rect 7300 13240 7328 13268
rect 6288 13212 7328 13240
rect 7644 13243 7702 13249
rect 6288 13172 6316 13212
rect 7644 13209 7656 13243
rect 7690 13240 7702 13243
rect 8202 13240 8208 13252
rect 7690 13212 8208 13240
rect 7690 13209 7702 13212
rect 7644 13203 7702 13209
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 10060 13240 10088 13416
rect 15396 13416 20628 13444
rect 10612 13348 11008 13376
rect 10612 13320 10640 13348
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 10980 13317 11008 13348
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 15396 13385 15424 13416
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 12952 13348 15393 13376
rect 12952 13336 12958 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 15838 13336 15844 13388
rect 15896 13336 15902 13388
rect 22572 13376 22600 13484
rect 25866 13472 25872 13484
rect 25924 13472 25930 13524
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 30561 13515 30619 13521
rect 30561 13512 30573 13515
rect 29420 13484 30573 13512
rect 29420 13472 29426 13484
rect 30561 13481 30573 13484
rect 30607 13481 30619 13515
rect 30561 13475 30619 13481
rect 15948 13348 22600 13376
rect 22741 13379 22799 13385
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11330 13308 11336 13320
rect 11103 13280 11336 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 10704 13240 10732 13271
rect 11330 13268 11336 13280
rect 11388 13308 11394 13320
rect 11882 13308 11888 13320
rect 11388 13280 11888 13308
rect 11388 13268 11394 13280
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 14458 13268 14464 13320
rect 14516 13308 14522 13320
rect 15194 13308 15200 13320
rect 14516 13280 15200 13308
rect 14516 13268 14522 13280
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15856 13308 15884 13336
rect 15335 13280 15884 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 10060 13212 10732 13240
rect 10873 13243 10931 13249
rect 10873 13209 10885 13243
rect 10919 13240 10931 13243
rect 11514 13240 11520 13252
rect 10919 13212 11520 13240
rect 10919 13209 10931 13212
rect 10873 13203 10931 13209
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 15948 13240 15976 13348
rect 22741 13345 22753 13379
rect 22787 13345 22799 13379
rect 22741 13339 22799 13345
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 22094 13308 22100 13320
rect 16172 13280 22100 13308
rect 16172 13268 16178 13280
rect 22094 13268 22100 13280
rect 22152 13308 22158 13320
rect 22756 13308 22784 13339
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 24949 13379 25007 13385
rect 24949 13376 24961 13379
rect 24728 13348 24961 13376
rect 24728 13336 24734 13348
rect 24949 13345 24961 13348
rect 24995 13345 25007 13379
rect 24949 13339 25007 13345
rect 22152 13280 22784 13308
rect 22152 13268 22158 13280
rect 23382 13268 23388 13320
rect 23440 13308 23446 13320
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 23440 13280 23489 13308
rect 23440 13268 23446 13280
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 25774 13268 25780 13320
rect 25832 13268 25838 13320
rect 14700 13212 15976 13240
rect 14700 13200 14706 13212
rect 18322 13200 18328 13252
rect 18380 13240 18386 13252
rect 18598 13240 18604 13252
rect 18380 13212 18604 13240
rect 18380 13200 18386 13212
rect 18598 13200 18604 13212
rect 18656 13200 18662 13252
rect 19426 13200 19432 13252
rect 19484 13240 19490 13252
rect 22370 13240 22376 13252
rect 19484 13212 22376 13240
rect 19484 13200 19490 13212
rect 22370 13200 22376 13212
rect 22428 13200 22434 13252
rect 22738 13200 22744 13252
rect 22796 13240 22802 13252
rect 30837 13243 30895 13249
rect 22796 13212 24808 13240
rect 22796 13200 22802 13212
rect 6104 13144 6316 13172
rect 6454 13132 6460 13184
rect 6512 13132 6518 13184
rect 7190 13132 7196 13184
rect 7248 13132 7254 13184
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 9950 13132 9956 13184
rect 10008 13132 10014 13184
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11330 13172 11336 13184
rect 11287 13144 11336 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11330 13132 11336 13144
rect 11388 13132 11394 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 15838 13172 15844 13184
rect 15252 13144 15844 13172
rect 15252 13132 15258 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 21450 13132 21456 13184
rect 21508 13172 21514 13184
rect 22097 13175 22155 13181
rect 22097 13172 22109 13175
rect 21508 13144 22109 13172
rect 21508 13132 21514 13144
rect 22097 13141 22109 13144
rect 22143 13141 22155 13175
rect 22388 13172 22416 13200
rect 24780 13184 24808 13212
rect 30837 13209 30849 13243
rect 30883 13240 30895 13243
rect 31294 13240 31300 13252
rect 30883 13212 31300 13240
rect 30883 13209 30895 13212
rect 30837 13203 30895 13209
rect 31294 13200 31300 13212
rect 31352 13200 31358 13252
rect 22465 13175 22523 13181
rect 22465 13172 22477 13175
rect 22388 13144 22477 13172
rect 22097 13135 22155 13141
rect 22465 13141 22477 13144
rect 22511 13141 22523 13175
rect 22465 13135 22523 13141
rect 22557 13175 22615 13181
rect 22557 13141 22569 13175
rect 22603 13172 22615 13175
rect 22925 13175 22983 13181
rect 22925 13172 22937 13175
rect 22603 13144 22937 13172
rect 22603 13141 22615 13144
rect 22557 13135 22615 13141
rect 22925 13141 22937 13144
rect 22971 13141 22983 13175
rect 22925 13135 22983 13141
rect 24394 13132 24400 13184
rect 24452 13132 24458 13184
rect 24762 13132 24768 13184
rect 24820 13132 24826 13184
rect 24857 13175 24915 13181
rect 24857 13141 24869 13175
rect 24903 13172 24915 13175
rect 25225 13175 25283 13181
rect 25225 13172 25237 13175
rect 24903 13144 25237 13172
rect 24903 13141 24915 13144
rect 24857 13135 24915 13141
rect 25225 13141 25237 13144
rect 25271 13141 25283 13175
rect 25225 13135 25283 13141
rect 1104 13082 31280 13104
rect 1104 13030 4922 13082
rect 4974 13030 4986 13082
rect 5038 13030 5050 13082
rect 5102 13030 5114 13082
rect 5166 13030 5178 13082
rect 5230 13030 5242 13082
rect 5294 13030 10922 13082
rect 10974 13030 10986 13082
rect 11038 13030 11050 13082
rect 11102 13030 11114 13082
rect 11166 13030 11178 13082
rect 11230 13030 11242 13082
rect 11294 13030 16922 13082
rect 16974 13030 16986 13082
rect 17038 13030 17050 13082
rect 17102 13030 17114 13082
rect 17166 13030 17178 13082
rect 17230 13030 17242 13082
rect 17294 13030 22922 13082
rect 22974 13030 22986 13082
rect 23038 13030 23050 13082
rect 23102 13030 23114 13082
rect 23166 13030 23178 13082
rect 23230 13030 23242 13082
rect 23294 13030 28922 13082
rect 28974 13030 28986 13082
rect 29038 13030 29050 13082
rect 29102 13030 29114 13082
rect 29166 13030 29178 13082
rect 29230 13030 29242 13082
rect 29294 13030 31280 13082
rect 1104 13008 31280 13030
rect 3329 12971 3387 12977
rect 3329 12937 3341 12971
rect 3375 12968 3387 12971
rect 3786 12968 3792 12980
rect 3375 12940 3792 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2038 12832 2044 12844
rect 1995 12804 2044 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2222 12841 2228 12844
rect 2216 12832 2228 12841
rect 2183 12804 2228 12832
rect 2216 12795 2228 12804
rect 2222 12792 2228 12795
rect 2280 12792 2286 12844
rect 3620 12841 3648 12940
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 3970 12928 3976 12980
rect 4028 12928 4034 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4706 12968 4712 12980
rect 4203 12940 4712 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5534 12928 5540 12980
rect 5592 12928 5598 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 6052 12940 6193 12968
rect 6052 12928 6058 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6365 12971 6423 12977
rect 6365 12937 6377 12971
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 7190 12968 7196 12980
rect 6779 12940 7196 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 3881 12903 3939 12909
rect 3881 12869 3893 12903
rect 3927 12900 3939 12903
rect 3988 12900 4016 12928
rect 5442 12900 5448 12912
rect 3927 12872 4016 12900
rect 4816 12872 5448 12900
rect 3927 12869 3939 12872
rect 3881 12863 3939 12869
rect 4816 12844 4844 12872
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 5552 12900 5580 12928
rect 6380 12900 6408 12931
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9030 12968 9036 12980
rect 7300 12940 9036 12968
rect 5552 12872 6408 12900
rect 6825 12903 6883 12909
rect 6825 12869 6837 12903
rect 6871 12900 6883 12903
rect 7006 12900 7012 12912
rect 6871 12872 7012 12900
rect 6871 12869 6883 12872
rect 6825 12863 6883 12869
rect 7006 12860 7012 12872
rect 7064 12900 7070 12912
rect 7300 12900 7328 12940
rect 9030 12928 9036 12940
rect 9088 12968 9094 12980
rect 9398 12968 9404 12980
rect 9088 12940 9404 12968
rect 9088 12928 9094 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 9950 12968 9956 12980
rect 9539 12940 9956 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10686 12928 10692 12980
rect 10744 12968 10750 12980
rect 10870 12968 10876 12980
rect 10744 12940 10876 12968
rect 10744 12928 10750 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 18598 12968 18604 12980
rect 17368 12940 18604 12968
rect 17368 12928 17374 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 19426 12928 19432 12980
rect 19484 12928 19490 12980
rect 21082 12928 21088 12980
rect 21140 12928 21146 12980
rect 21266 12928 21272 12980
rect 21324 12928 21330 12980
rect 21358 12928 21364 12980
rect 21416 12928 21422 12980
rect 21637 12971 21695 12977
rect 21637 12937 21649 12971
rect 21683 12968 21695 12971
rect 23201 12971 23259 12977
rect 21683 12940 22094 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 7064 12872 7328 12900
rect 7064 12860 7070 12872
rect 7374 12860 7380 12912
rect 7432 12900 7438 12912
rect 7926 12900 7932 12912
rect 7432 12872 7932 12900
rect 7432 12860 7438 12872
rect 7926 12860 7932 12872
rect 7984 12860 7990 12912
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 8803 12872 10456 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12801 3663 12835
rect 3605 12795 3663 12801
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4019 12804 4752 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 3804 12764 3832 12795
rect 4522 12764 4528 12776
rect 3804 12736 4528 12764
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4724 12628 4752 12804
rect 4798 12792 4804 12844
rect 4856 12792 4862 12844
rect 5068 12835 5126 12841
rect 5068 12801 5080 12835
rect 5114 12832 5126 12835
rect 5350 12832 5356 12844
rect 5114 12804 5356 12832
rect 5114 12801 5126 12804
rect 5068 12795 5126 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 10428 12841 10456 12872
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10502 12832 10508 12844
rect 10459 12804 10508 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10502 12792 10508 12804
rect 10560 12792 10566 12844
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 6822 12764 6828 12776
rect 6696 12736 6828 12764
rect 6696 12724 6702 12736
rect 6822 12724 6828 12736
rect 6880 12764 6886 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6880 12736 6929 12764
rect 6880 12724 6886 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 10704 12764 10732 12928
rect 10962 12860 10968 12912
rect 11020 12900 11026 12912
rect 11241 12903 11299 12909
rect 11241 12900 11253 12903
rect 11020 12872 11253 12900
rect 11020 12860 11026 12872
rect 11241 12869 11253 12872
rect 11287 12900 11299 12903
rect 11606 12900 11612 12912
rect 11287 12872 11612 12900
rect 11287 12869 11299 12872
rect 11241 12863 11299 12869
rect 11606 12860 11612 12872
rect 11664 12900 11670 12912
rect 14090 12900 14096 12912
rect 11664 12872 14096 12900
rect 11664 12860 11670 12872
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 20993 12903 21051 12909
rect 19076 12872 20852 12900
rect 19076 12844 19104 12872
rect 17034 12792 17040 12844
rect 17092 12792 17098 12844
rect 19058 12792 19064 12844
rect 19116 12792 19122 12844
rect 19521 12835 19579 12841
rect 19521 12801 19533 12835
rect 19567 12832 19579 12835
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19567 12804 19993 12832
rect 19567 12801 19579 12804
rect 19521 12795 19579 12801
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20824 12841 20852 12872
rect 20993 12869 21005 12903
rect 21039 12900 21051 12903
rect 21100 12900 21128 12928
rect 21039 12872 21128 12900
rect 21284 12900 21312 12928
rect 22066 12909 22094 12940
rect 23201 12937 23213 12971
rect 23247 12968 23259 12971
rect 23382 12968 23388 12980
rect 23247 12940 23388 12968
rect 23247 12937 23259 12940
rect 23201 12931 23259 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 23753 12971 23811 12977
rect 23753 12937 23765 12971
rect 23799 12937 23811 12971
rect 23753 12931 23811 12937
rect 22066 12903 22124 12909
rect 21284 12872 21864 12900
rect 21039 12869 21051 12872
rect 20993 12863 21051 12869
rect 21836 12844 21864 12872
rect 22066 12869 22078 12903
rect 22112 12869 22124 12903
rect 23474 12900 23480 12912
rect 22066 12863 22124 12869
rect 23216 12872 23480 12900
rect 23216 12844 23244 12872
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 23768 12900 23796 12931
rect 24394 12928 24400 12980
rect 24452 12928 24458 12980
rect 25222 12928 25228 12980
rect 25280 12968 25286 12980
rect 25774 12968 25780 12980
rect 25280 12940 25780 12968
rect 25280 12928 25286 12940
rect 25774 12928 25780 12940
rect 25832 12928 25838 12980
rect 26418 12928 26424 12980
rect 26476 12928 26482 12980
rect 29362 12928 29368 12980
rect 29420 12928 29426 12980
rect 24090 12903 24148 12909
rect 24090 12900 24102 12903
rect 23768 12872 24102 12900
rect 24090 12869 24102 12872
rect 24136 12869 24148 12903
rect 24090 12863 24148 12869
rect 20717 12835 20775 12841
rect 20717 12832 20729 12835
rect 20404 12804 20729 12832
rect 20404 12792 20410 12804
rect 20717 12801 20729 12804
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 20810 12835 20868 12841
rect 20810 12801 20822 12835
rect 20856 12801 20868 12835
rect 20810 12795 20868 12801
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12801 21143 12835
rect 21085 12795 21143 12801
rect 9631 12736 10732 12764
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11422 12764 11428 12776
rect 11204 12736 11428 12764
rect 11204 12724 11210 12736
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 17126 12724 17132 12776
rect 17184 12724 17190 12776
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12764 17371 12767
rect 17494 12764 17500 12776
rect 17359 12736 17500 12764
rect 17359 12733 17371 12736
rect 17313 12727 17371 12733
rect 17494 12724 17500 12736
rect 17552 12764 17558 12776
rect 17770 12764 17776 12776
rect 17552 12736 17776 12764
rect 17552 12724 17558 12736
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18138 12724 18144 12776
rect 18196 12724 18202 12776
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19794 12764 19800 12776
rect 19383 12736 19800 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19794 12724 19800 12736
rect 19852 12724 19858 12776
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 21100 12764 21128 12795
rect 21174 12792 21180 12844
rect 21232 12841 21238 12844
rect 21232 12832 21240 12841
rect 21232 12804 21277 12832
rect 21232 12795 21240 12804
rect 21232 12792 21238 12795
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 21818 12792 21824 12844
rect 21876 12792 21882 12844
rect 23198 12792 23204 12844
rect 23256 12792 23262 12844
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 23569 12835 23627 12841
rect 23569 12801 23581 12835
rect 23615 12832 23627 12835
rect 24412 12832 24440 12928
rect 24762 12860 24768 12912
rect 24820 12900 24826 12912
rect 25685 12903 25743 12909
rect 25685 12900 25697 12903
rect 24820 12872 25697 12900
rect 24820 12860 24826 12872
rect 25685 12869 25697 12872
rect 25731 12900 25743 12903
rect 26436 12900 26464 12928
rect 25731 12872 26464 12900
rect 25731 12869 25743 12872
rect 25685 12863 25743 12869
rect 23615 12804 24440 12832
rect 25777 12835 25835 12841
rect 23615 12801 23627 12804
rect 23569 12795 23627 12801
rect 25777 12801 25789 12835
rect 25823 12832 25835 12835
rect 26145 12835 26203 12841
rect 26145 12832 26157 12835
rect 25823 12804 26157 12832
rect 25823 12801 25835 12804
rect 25777 12795 25835 12801
rect 26145 12801 26157 12804
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 28629 12835 28687 12841
rect 28629 12801 28641 12835
rect 28675 12832 28687 12835
rect 29380 12832 29408 12928
rect 28675 12804 29408 12832
rect 28675 12801 28687 12804
rect 28629 12795 28687 12801
rect 20680 12736 21128 12764
rect 20680 12724 20686 12736
rect 6454 12656 6460 12708
rect 6512 12696 6518 12708
rect 6512 12668 11468 12696
rect 6512 12656 6518 12668
rect 11440 12640 11468 12668
rect 19702 12656 19708 12708
rect 19760 12696 19766 12708
rect 23308 12696 23336 12795
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23532 12736 23857 12764
rect 23532 12724 23538 12736
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 23845 12727 23903 12733
rect 25866 12724 25872 12776
rect 25924 12724 25930 12776
rect 26694 12724 26700 12776
rect 26752 12724 26758 12776
rect 28074 12724 28080 12776
rect 28132 12724 28138 12776
rect 19760 12668 21864 12696
rect 23308 12668 23796 12696
rect 19760 12656 19766 12668
rect 5534 12628 5540 12640
rect 4724 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 9033 12631 9091 12637
rect 9033 12628 9045 12631
rect 8904 12600 9045 12628
rect 8904 12588 8910 12600
rect 9033 12597 9045 12600
rect 9079 12597 9091 12631
rect 9033 12591 9091 12597
rect 11422 12588 11428 12640
rect 11480 12588 11486 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 11882 12628 11888 12640
rect 11756 12600 11888 12628
rect 11756 12588 11762 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 13722 12588 13728 12640
rect 13780 12588 13786 12640
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 17586 12588 17592 12640
rect 17644 12588 17650 12640
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 18690 12628 18696 12640
rect 18463 12600 18696 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20714 12628 20720 12640
rect 19935 12600 20720 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21836 12628 21864 12668
rect 22738 12628 22744 12640
rect 21836 12600 22744 12628
rect 22738 12588 22744 12600
rect 22796 12628 22802 12640
rect 23106 12628 23112 12640
rect 22796 12600 23112 12628
rect 22796 12588 22802 12600
rect 23106 12588 23112 12600
rect 23164 12588 23170 12640
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 23658 12628 23664 12640
rect 23523 12600 23664 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 23658 12588 23664 12600
rect 23716 12588 23722 12640
rect 23768 12628 23796 12668
rect 25317 12631 25375 12637
rect 25317 12628 25329 12631
rect 23768 12600 25329 12628
rect 25317 12597 25329 12600
rect 25363 12597 25375 12631
rect 25317 12591 25375 12597
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 27433 12631 27491 12637
rect 27433 12628 27445 12631
rect 26476 12600 27445 12628
rect 26476 12588 26482 12600
rect 27433 12597 27445 12600
rect 27479 12597 27491 12631
rect 27433 12591 27491 12597
rect 28537 12631 28595 12637
rect 28537 12597 28549 12631
rect 28583 12628 28595 12631
rect 28626 12628 28632 12640
rect 28583 12600 28632 12628
rect 28583 12597 28595 12600
rect 28537 12591 28595 12597
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 1104 12538 31280 12560
rect 1104 12486 4182 12538
rect 4234 12486 4246 12538
rect 4298 12486 4310 12538
rect 4362 12486 4374 12538
rect 4426 12486 4438 12538
rect 4490 12486 4502 12538
rect 4554 12486 10182 12538
rect 10234 12486 10246 12538
rect 10298 12486 10310 12538
rect 10362 12486 10374 12538
rect 10426 12486 10438 12538
rect 10490 12486 10502 12538
rect 10554 12486 16182 12538
rect 16234 12486 16246 12538
rect 16298 12486 16310 12538
rect 16362 12486 16374 12538
rect 16426 12486 16438 12538
rect 16490 12486 16502 12538
rect 16554 12486 22182 12538
rect 22234 12486 22246 12538
rect 22298 12486 22310 12538
rect 22362 12486 22374 12538
rect 22426 12486 22438 12538
rect 22490 12486 22502 12538
rect 22554 12486 28182 12538
rect 28234 12486 28246 12538
rect 28298 12486 28310 12538
rect 28362 12486 28374 12538
rect 28426 12486 28438 12538
rect 28490 12486 28502 12538
rect 28554 12486 31280 12538
rect 1104 12464 31280 12486
rect 5442 12424 5448 12436
rect 5092 12396 5448 12424
rect 5092 12297 5120 12396
rect 5442 12384 5448 12396
rect 5500 12424 5506 12436
rect 7926 12424 7932 12436
rect 5500 12396 7932 12424
rect 5500 12384 5506 12396
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8202 12384 8208 12436
rect 8260 12384 8266 12436
rect 10321 12427 10379 12433
rect 10321 12393 10333 12427
rect 10367 12424 10379 12427
rect 10594 12424 10600 12436
rect 10367 12396 10600 12424
rect 10367 12393 10379 12396
rect 10321 12387 10379 12393
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 10686 12384 10692 12436
rect 10744 12384 10750 12436
rect 11330 12424 11336 12436
rect 11164 12396 11336 12424
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 6457 12359 6515 12365
rect 6457 12356 6469 12359
rect 6236 12328 6469 12356
rect 6236 12316 6242 12328
rect 6457 12325 6469 12328
rect 6503 12356 6515 12359
rect 8938 12356 8944 12368
rect 6503 12328 7972 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 5077 12291 5135 12297
rect 5077 12257 5089 12291
rect 5123 12257 5135 12291
rect 5077 12251 5135 12257
rect 6822 12248 6828 12300
rect 6880 12248 6886 12300
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 7944 12297 7972 12328
rect 8404 12328 8944 12356
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 6840 12220 6868 12248
rect 7116 12220 7144 12251
rect 8404 12229 8432 12328
rect 8938 12316 8944 12328
rect 8996 12316 9002 12368
rect 10502 12316 10508 12368
rect 10560 12356 10566 12368
rect 10704 12356 10732 12384
rect 10560 12328 10732 12356
rect 10560 12316 10566 12328
rect 11164 12288 11192 12396
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17092 12396 17509 12424
rect 17092 12384 17098 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 19061 12427 19119 12433
rect 19061 12393 19073 12427
rect 19107 12424 19119 12427
rect 19107 12396 20576 12424
rect 19107 12393 19119 12396
rect 19061 12387 19119 12393
rect 11241 12359 11299 12365
rect 11241 12325 11253 12359
rect 11287 12356 11299 12359
rect 11701 12359 11759 12365
rect 11287 12328 11468 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 11440 12297 11468 12328
rect 11701 12325 11713 12359
rect 11747 12356 11759 12359
rect 13446 12356 13452 12368
rect 11747 12328 12434 12356
rect 11747 12325 11759 12328
rect 11701 12319 11759 12325
rect 10612 12260 11192 12288
rect 11425 12291 11483 12297
rect 6840 12192 7144 12220
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8846 12220 8852 12232
rect 8619 12192 8852 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8846 12180 8852 12192
rect 8904 12180 8910 12232
rect 10612 12229 10640 12260
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 12406 12288 12434 12328
rect 13280 12328 13452 12356
rect 13280 12297 13308 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 13265 12291 13323 12297
rect 12406 12260 12480 12288
rect 11425 12251 11483 12257
rect 8941 12223 8999 12229
rect 8941 12189 8953 12223
rect 8987 12220 8999 12223
rect 10597 12223 10655 12229
rect 8987 12192 9674 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 5344 12155 5402 12161
rect 5344 12121 5356 12155
rect 5390 12152 5402 12155
rect 5534 12152 5540 12164
rect 5390 12124 5540 12152
rect 5390 12121 5402 12124
rect 5344 12115 5402 12121
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 9186 12155 9244 12161
rect 9186 12152 9198 12155
rect 8772 12124 9198 12152
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5442 12084 5448 12096
rect 4764 12056 5448 12084
rect 4764 12044 4770 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6546 12044 6552 12096
rect 6604 12044 6610 12096
rect 8772 12093 8800 12124
rect 9186 12121 9198 12124
rect 9232 12121 9244 12155
rect 9186 12115 9244 12121
rect 9646 12096 9674 12192
rect 10597 12189 10609 12223
rect 10643 12189 10655 12223
rect 10597 12183 10655 12189
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10796 12192 10977 12220
rect 10410 12112 10416 12164
rect 10468 12152 10474 12164
rect 10796 12152 10824 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11062 12223 11120 12229
rect 11062 12189 11074 12223
rect 11108 12220 11120 12223
rect 11333 12223 11391 12229
rect 11108 12192 11192 12220
rect 11108 12189 11120 12192
rect 11062 12183 11120 12189
rect 10468 12124 10824 12152
rect 10873 12155 10931 12161
rect 10468 12112 10474 12124
rect 10873 12121 10885 12155
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7377 12087 7435 12093
rect 7377 12084 7389 12087
rect 6963 12056 7389 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7377 12053 7389 12056
rect 7423 12053 7435 12087
rect 7377 12047 7435 12053
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12053 8815 12087
rect 9646 12056 9680 12096
rect 8757 12047 8815 12053
rect 9674 12044 9680 12056
rect 9732 12084 9738 12096
rect 10778 12084 10784 12096
rect 9732 12056 10784 12084
rect 9732 12044 9738 12056
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 10888 12084 10916 12115
rect 11054 12084 11060 12096
rect 10888 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11164 12084 11192 12192
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 12066 12220 12072 12232
rect 11379 12192 12072 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12250 12180 12256 12232
rect 12308 12180 12314 12232
rect 12452 12229 12480 12260
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 13722 12288 13728 12300
rect 13403 12260 13728 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17402 12288 17408 12300
rect 17359 12260 17408 12288
rect 17359 12257 17371 12260
rect 17313 12251 17371 12257
rect 17402 12248 17408 12260
rect 17460 12288 17466 12300
rect 17678 12288 17684 12300
rect 17460 12260 17684 12288
rect 17460 12248 17466 12260
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 18414 12248 18420 12300
rect 18472 12248 18478 12300
rect 20548 12288 20576 12396
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 23566 12424 23572 12436
rect 21784 12396 23572 12424
rect 21784 12384 21790 12396
rect 23566 12384 23572 12396
rect 23624 12384 23630 12436
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 24026 12424 24032 12436
rect 23716 12396 24032 12424
rect 23716 12384 23722 12396
rect 24026 12384 24032 12396
rect 24084 12384 24090 12436
rect 24210 12384 24216 12436
rect 24268 12384 24274 12436
rect 25777 12427 25835 12433
rect 25777 12424 25789 12427
rect 24412 12396 25789 12424
rect 23198 12316 23204 12368
rect 23256 12316 23262 12368
rect 24412 12356 24440 12396
rect 25777 12393 25789 12396
rect 25823 12424 25835 12427
rect 26694 12424 26700 12436
rect 25823 12396 26700 12424
rect 25823 12393 25835 12396
rect 25777 12387 25835 12393
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 29089 12427 29147 12433
rect 29089 12393 29101 12427
rect 29135 12424 29147 12427
rect 30650 12424 30656 12436
rect 29135 12396 30656 12424
rect 29135 12393 29147 12396
rect 29089 12387 29147 12393
rect 30650 12384 30656 12396
rect 30708 12384 30714 12436
rect 23860 12328 24440 12356
rect 20548 12260 21220 12288
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12220 12679 12223
rect 15378 12220 15384 12232
rect 12667 12192 15384 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12220 17095 12223
rect 17586 12220 17592 12232
rect 17083 12192 17592 12220
rect 17083 12189 17095 12192
rect 17037 12183 17095 12189
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 12345 12155 12403 12161
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 14182 12152 14188 12164
rect 12391 12124 14188 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 18064 12096 18092 12183
rect 18432 12152 18460 12248
rect 18690 12180 18696 12232
rect 18748 12180 18754 12232
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19291 12192 19656 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19334 12152 19340 12164
rect 18432 12124 19340 12152
rect 19334 12112 19340 12124
rect 19392 12112 19398 12164
rect 19512 12155 19570 12161
rect 19512 12121 19524 12155
rect 19558 12121 19570 12155
rect 19628 12152 19656 12192
rect 20898 12180 20904 12232
rect 20956 12180 20962 12232
rect 21192 12229 21220 12260
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21450 12180 21456 12232
rect 21508 12180 21514 12232
rect 22945 12223 23003 12229
rect 22945 12220 22957 12223
rect 22940 12189 22957 12220
rect 22991 12189 23003 12223
rect 23216 12220 23244 12316
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 23216 12192 23305 12220
rect 22940 12183 23003 12189
rect 23293 12189 23305 12192
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 21468 12152 21496 12180
rect 21726 12161 21732 12164
rect 19628 12124 21496 12152
rect 19512 12115 19570 12121
rect 21720 12115 21732 12161
rect 11606 12084 11612 12096
rect 11164 12056 11612 12084
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 12066 12044 12072 12096
rect 12124 12044 12130 12096
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 13449 12087 13507 12093
rect 13449 12084 13461 12087
rect 12768 12056 13461 12084
rect 12768 12044 12774 12056
rect 13449 12053 13461 12056
rect 13495 12053 13507 12087
rect 13449 12047 13507 12053
rect 13814 12044 13820 12096
rect 13872 12044 13878 12096
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17862 12084 17868 12096
rect 17184 12056 17868 12084
rect 17184 12044 17190 12056
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 18046 12044 18052 12096
rect 18104 12044 18110 12096
rect 18601 12087 18659 12093
rect 18601 12053 18613 12087
rect 18647 12084 18659 12087
rect 19426 12084 19432 12096
rect 18647 12056 19432 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 19536 12084 19564 12115
rect 21726 12112 21732 12115
rect 21784 12112 21790 12164
rect 22940 12152 22968 12183
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 23569 12223 23627 12229
rect 23569 12220 23581 12223
rect 23492 12192 23581 12220
rect 22940 12124 23060 12152
rect 20717 12087 20775 12093
rect 20717 12084 20729 12087
rect 19536 12056 20729 12084
rect 20717 12053 20729 12056
rect 20763 12053 20775 12087
rect 20717 12047 20775 12053
rect 20990 12044 20996 12096
rect 21048 12044 21054 12096
rect 22833 12087 22891 12093
rect 22833 12053 22845 12087
rect 22879 12084 22891 12087
rect 23032 12084 23060 12124
rect 23106 12112 23112 12164
rect 23164 12112 23170 12164
rect 23201 12155 23259 12161
rect 23201 12121 23213 12155
rect 23247 12152 23259 12155
rect 23400 12152 23428 12180
rect 23247 12124 23428 12152
rect 23247 12121 23259 12124
rect 23201 12115 23259 12121
rect 23382 12084 23388 12096
rect 22879 12056 23388 12084
rect 22879 12053 22891 12056
rect 22833 12047 22891 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 23492 12093 23520 12192
rect 23569 12189 23581 12192
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 23717 12223 23775 12229
rect 23717 12189 23729 12223
rect 23763 12220 23775 12223
rect 23860 12220 23888 12328
rect 26234 12248 26240 12300
rect 26292 12288 26298 12300
rect 26292 12260 27016 12288
rect 26292 12248 26298 12260
rect 23763 12192 23888 12220
rect 23937 12223 23995 12229
rect 23763 12189 23775 12192
rect 23717 12183 23775 12189
rect 23937 12189 23949 12223
rect 23983 12189 23995 12223
rect 23937 12183 23995 12189
rect 24075 12223 24133 12229
rect 24075 12189 24087 12223
rect 24121 12220 24133 12223
rect 24302 12220 24308 12232
rect 24121 12192 24308 12220
rect 24121 12189 24133 12192
rect 24075 12183 24133 12189
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12121 23903 12155
rect 23845 12115 23903 12121
rect 23477 12087 23535 12093
rect 23477 12053 23489 12087
rect 23523 12053 23535 12087
rect 23477 12047 23535 12053
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23860 12084 23888 12115
rect 23624 12056 23888 12084
rect 23952 12084 23980 12183
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12220 24455 12223
rect 24486 12220 24492 12232
rect 24443 12192 24492 12220
rect 24443 12189 24455 12192
rect 24397 12183 24455 12189
rect 24486 12180 24492 12192
rect 24544 12220 24550 12232
rect 26252 12220 26280 12248
rect 26988 12232 27016 12260
rect 24544 12192 26280 12220
rect 24544 12180 24550 12192
rect 26418 12180 26424 12232
rect 26476 12180 26482 12232
rect 26513 12223 26571 12229
rect 26513 12189 26525 12223
rect 26559 12220 26571 12223
rect 26602 12220 26608 12232
rect 26559 12192 26608 12220
rect 26559 12189 26571 12192
rect 26513 12183 26571 12189
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 26694 12180 26700 12232
rect 26752 12180 26758 12232
rect 26970 12180 26976 12232
rect 27028 12220 27034 12232
rect 27341 12223 27399 12229
rect 27341 12220 27353 12223
rect 27028 12192 27353 12220
rect 27028 12180 27034 12192
rect 27341 12189 27353 12192
rect 27387 12189 27399 12223
rect 27341 12183 27399 12189
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 24642 12155 24700 12161
rect 24642 12152 24654 12155
rect 24268 12124 24654 12152
rect 24268 12112 24274 12124
rect 24642 12121 24654 12124
rect 24688 12121 24700 12155
rect 24642 12115 24700 12121
rect 26142 12112 26148 12164
rect 26200 12152 26206 12164
rect 26712 12152 26740 12180
rect 26200 12124 26740 12152
rect 26200 12112 26206 12124
rect 27614 12112 27620 12164
rect 27672 12112 27678 12164
rect 28626 12112 28632 12164
rect 28684 12112 28690 12164
rect 25222 12084 25228 12096
rect 23952 12056 25228 12084
rect 23624 12044 23630 12056
rect 25222 12044 25228 12056
rect 25280 12044 25286 12096
rect 26878 12044 26884 12096
rect 26936 12044 26942 12096
rect 1104 11994 31280 12016
rect 1104 11942 4922 11994
rect 4974 11942 4986 11994
rect 5038 11942 5050 11994
rect 5102 11942 5114 11994
rect 5166 11942 5178 11994
rect 5230 11942 5242 11994
rect 5294 11942 10922 11994
rect 10974 11942 10986 11994
rect 11038 11942 11050 11994
rect 11102 11942 11114 11994
rect 11166 11942 11178 11994
rect 11230 11942 11242 11994
rect 11294 11942 16922 11994
rect 16974 11942 16986 11994
rect 17038 11942 17050 11994
rect 17102 11942 17114 11994
rect 17166 11942 17178 11994
rect 17230 11942 17242 11994
rect 17294 11942 22922 11994
rect 22974 11942 22986 11994
rect 23038 11942 23050 11994
rect 23102 11942 23114 11994
rect 23166 11942 23178 11994
rect 23230 11942 23242 11994
rect 23294 11942 28922 11994
rect 28974 11942 28986 11994
rect 29038 11942 29050 11994
rect 29102 11942 29114 11994
rect 29166 11942 29178 11994
rect 29230 11942 29242 11994
rect 29294 11942 31280 11994
rect 1104 11920 31280 11942
rect 5534 11840 5540 11892
rect 5592 11840 5598 11892
rect 6546 11840 6552 11892
rect 6604 11840 6610 11892
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 992 11716 1409 11744
rect 992 11704 998 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 3973 11747 4031 11753
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4798 11744 4804 11756
rect 4019 11716 4804 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 1780 11676 1808 11707
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 6564 11744 6592 11840
rect 5767 11716 6592 11744
rect 8573 11747 8631 11753
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8864 11744 8892 11843
rect 10502 11840 10508 11892
rect 10560 11880 10566 11892
rect 10870 11880 10876 11892
rect 10560 11852 10876 11880
rect 10560 11840 10566 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 15378 11840 15384 11892
rect 15436 11840 15442 11892
rect 16666 11880 16672 11892
rect 16316 11852 16672 11880
rect 8619 11716 8892 11744
rect 9217 11747 9275 11753
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9582 11744 9588 11756
rect 9263 11716 9588 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9674 11704 9680 11756
rect 9732 11704 9738 11756
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 9944 11747 10002 11753
rect 9944 11713 9956 11747
rect 9990 11744 10002 11747
rect 9990 11716 10732 11744
rect 9990 11713 10002 11716
rect 9944 11707 10002 11713
rect 9309 11679 9367 11685
rect 1780 11648 8892 11676
rect 3786 11500 3792 11552
rect 3844 11500 3850 11552
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 8864 11540 8892 11648
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9493 11679 9551 11685
rect 9493 11645 9505 11679
rect 9539 11676 9551 11679
rect 9784 11676 9812 11704
rect 9539 11648 9812 11676
rect 9539 11645 9551 11648
rect 9493 11639 9551 11645
rect 9324 11608 9352 11639
rect 9674 11608 9680 11620
rect 9324 11580 9680 11608
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 10704 11608 10732 11716
rect 10888 11676 10916 11840
rect 11330 11704 11336 11756
rect 11388 11704 11394 11756
rect 12084 11753 12112 11840
rect 13832 11812 13860 11840
rect 13832 11784 15700 11812
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 13837 11747 13895 11753
rect 13837 11713 13849 11747
rect 13883 11744 13895 11747
rect 13883 11716 14044 11744
rect 13883 11713 13895 11716
rect 13837 11707 13895 11713
rect 14016 11676 14044 11716
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14734 11704 14740 11756
rect 14792 11704 14798 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15672 11753 15700 11784
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14884 11716 15025 11744
rect 14884 11704 14890 11716
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 14921 11679 14979 11685
rect 14921 11676 14933 11679
rect 10888 11648 12434 11676
rect 14016 11648 14136 11676
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10704 11580 11161 11608
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 11149 11571 11207 11577
rect 11882 11568 11888 11620
rect 11940 11608 11946 11620
rect 12250 11608 12256 11620
rect 11940 11580 12256 11608
rect 11940 11568 11946 11580
rect 12250 11568 12256 11580
rect 12308 11568 12314 11620
rect 12406 11608 12434 11648
rect 14108 11620 14136 11648
rect 14200 11648 14933 11676
rect 12894 11608 12900 11620
rect 12406 11580 12900 11608
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 14090 11568 14096 11620
rect 14148 11568 14154 11620
rect 9950 11540 9956 11552
rect 8864 11512 9956 11540
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 11057 11543 11115 11549
rect 11057 11540 11069 11543
rect 10468 11512 11069 11540
rect 10468 11500 10474 11512
rect 11057 11509 11069 11512
rect 11103 11540 11115 11543
rect 11790 11540 11796 11552
rect 11103 11512 11796 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12621 11543 12679 11549
rect 12621 11540 12633 11543
rect 12584 11512 12633 11540
rect 12584 11500 12590 11512
rect 12621 11509 12633 11512
rect 12667 11509 12679 11543
rect 12621 11503 12679 11509
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11540 12771 11543
rect 13170 11540 13176 11552
rect 12759 11512 13176 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 13170 11500 13176 11512
rect 13228 11540 13234 11552
rect 14200 11540 14228 11648
rect 14921 11645 14933 11648
rect 14967 11645 14979 11679
rect 15212 11676 15240 11707
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 16316 11753 16344 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 18138 11880 18144 11892
rect 18095 11852 18144 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18969 11883 19027 11889
rect 18969 11849 18981 11883
rect 19015 11880 19027 11883
rect 19058 11880 19064 11892
rect 19015 11852 19064 11880
rect 19015 11849 19027 11852
rect 18969 11843 19027 11849
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 21450 11840 21456 11892
rect 21508 11840 21514 11892
rect 21637 11883 21695 11889
rect 21637 11849 21649 11883
rect 21683 11880 21695 11883
rect 21726 11880 21732 11892
rect 21683 11852 21732 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 23474 11880 23480 11892
rect 22664 11852 23480 11880
rect 16758 11812 16764 11824
rect 16684 11784 16764 11812
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11713 16359 11747
rect 16574 11744 16580 11756
rect 16301 11707 16359 11713
rect 16408 11716 16580 11744
rect 15286 11676 15292 11688
rect 15212 11648 15292 11676
rect 14921 11639 14979 11645
rect 15286 11636 15292 11648
rect 15344 11676 15350 11688
rect 16040 11676 16068 11704
rect 15344 11648 16068 11676
rect 16224 11676 16252 11707
rect 16408 11676 16436 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16684 11753 16712 11784
rect 16758 11772 16764 11784
rect 16816 11812 16822 11824
rect 21468 11812 21496 11840
rect 16816 11784 21496 11812
rect 16816 11772 16822 11784
rect 20364 11756 20392 11784
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 22664 11821 22692 11852
rect 23474 11840 23480 11852
rect 23532 11880 23538 11892
rect 24486 11880 24492 11892
rect 23532 11852 24492 11880
rect 23532 11840 23538 11852
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 26053 11883 26111 11889
rect 26053 11849 26065 11883
rect 26099 11849 26111 11883
rect 26053 11843 26111 11849
rect 22649 11815 22707 11821
rect 22649 11812 22661 11815
rect 21968 11784 22661 11812
rect 21968 11772 21974 11784
rect 22649 11781 22661 11784
rect 22695 11781 22707 11815
rect 22649 11775 22707 11781
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 16925 11747 16983 11753
rect 16925 11744 16937 11747
rect 16669 11707 16727 11713
rect 16776 11716 16937 11744
rect 16776 11676 16804 11716
rect 16925 11713 16937 11716
rect 16971 11713 16983 11747
rect 18046 11744 18052 11756
rect 16925 11707 16983 11713
rect 17880 11716 18052 11744
rect 16224 11648 16436 11676
rect 16500 11648 16804 11676
rect 15344 11636 15350 11648
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 16500 11617 16528 11648
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 14332 11580 15485 11608
rect 14332 11568 14338 11580
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 15473 11571 15531 11577
rect 16485 11611 16543 11617
rect 16485 11577 16497 11611
rect 16531 11577 16543 11611
rect 16485 11571 16543 11577
rect 13228 11512 14228 11540
rect 13228 11500 13234 11512
rect 16022 11500 16028 11552
rect 16080 11500 16086 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17880 11540 17908 11716
rect 18046 11704 18052 11716
rect 18104 11744 18110 11756
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 18104 11716 18153 11744
rect 18104 11704 18110 11716
rect 18141 11713 18153 11716
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18230 11704 18236 11756
rect 18288 11704 18294 11756
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11744 18567 11747
rect 18598 11744 18604 11756
rect 18555 11716 18604 11744
rect 18555 11713 18567 11716
rect 18509 11707 18567 11713
rect 18248 11676 18276 11704
rect 18432 11676 18460 11707
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 20093 11747 20151 11753
rect 20093 11713 20105 11747
rect 20139 11744 20151 11747
rect 20139 11716 20300 11744
rect 20139 11713 20151 11716
rect 20093 11707 20151 11713
rect 18248 11648 18460 11676
rect 20272 11676 20300 11716
rect 20346 11704 20352 11756
rect 20404 11704 20410 11756
rect 20990 11704 20996 11756
rect 21048 11704 21054 11756
rect 21450 11704 21456 11756
rect 21508 11704 21514 11756
rect 21542 11704 21548 11756
rect 21600 11744 21606 11756
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21600 11716 21833 11744
rect 21600 11704 21606 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 23382 11704 23388 11756
rect 23440 11704 23446 11756
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11744 25835 11747
rect 26068 11744 26096 11843
rect 26418 11840 26424 11892
rect 26476 11880 26482 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26476 11852 26525 11880
rect 26476 11840 26482 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 26513 11843 26571 11849
rect 28074 11840 28080 11892
rect 28132 11880 28138 11892
rect 28353 11883 28411 11889
rect 28353 11880 28365 11883
rect 28132 11852 28365 11880
rect 28132 11840 28138 11852
rect 28353 11849 28365 11852
rect 28399 11849 28411 11883
rect 28353 11843 28411 11849
rect 25823 11716 26096 11744
rect 25823 11713 25835 11716
rect 25777 11707 25835 11713
rect 26418 11704 26424 11756
rect 26476 11704 26482 11756
rect 27229 11747 27287 11753
rect 27229 11744 27241 11747
rect 26528 11716 27241 11744
rect 21008 11676 21036 11704
rect 20272 11648 21036 11676
rect 20438 11568 20444 11620
rect 20496 11568 20502 11620
rect 25961 11611 26019 11617
rect 25961 11577 25973 11611
rect 26007 11608 26019 11611
rect 26528 11608 26556 11716
rect 27229 11713 27241 11716
rect 27275 11713 27287 11747
rect 27229 11707 27287 11713
rect 30650 11704 30656 11756
rect 30708 11704 30714 11756
rect 26697 11679 26755 11685
rect 26697 11645 26709 11679
rect 26743 11645 26755 11679
rect 26697 11639 26755 11645
rect 26007 11580 26556 11608
rect 26007 11577 26019 11580
rect 25961 11571 26019 11577
rect 17368 11512 17908 11540
rect 18693 11543 18751 11549
rect 17368 11500 17374 11512
rect 18693 11509 18705 11543
rect 18739 11540 18751 11543
rect 20456 11540 20484 11568
rect 18739 11512 20484 11540
rect 18739 11509 18751 11512
rect 18693 11503 18751 11509
rect 22646 11500 22652 11552
rect 22704 11540 22710 11552
rect 22833 11543 22891 11549
rect 22833 11540 22845 11543
rect 22704 11512 22845 11540
rect 22704 11500 22710 11512
rect 22833 11509 22845 11512
rect 22879 11509 22891 11543
rect 22833 11503 22891 11509
rect 26326 11500 26332 11552
rect 26384 11540 26390 11552
rect 26510 11540 26516 11552
rect 26384 11512 26516 11540
rect 26384 11500 26390 11512
rect 26510 11500 26516 11512
rect 26568 11540 26574 11552
rect 26712 11540 26740 11639
rect 26970 11636 26976 11688
rect 27028 11636 27034 11688
rect 29089 11679 29147 11685
rect 29089 11645 29101 11679
rect 29135 11676 29147 11679
rect 30668 11676 30696 11704
rect 29135 11648 30696 11676
rect 29135 11645 29147 11648
rect 29089 11639 29147 11645
rect 26568 11512 26740 11540
rect 26568 11500 26574 11512
rect 27706 11500 27712 11552
rect 27764 11540 27770 11552
rect 28445 11543 28503 11549
rect 28445 11540 28457 11543
rect 27764 11512 28457 11540
rect 27764 11500 27770 11512
rect 28445 11509 28457 11512
rect 28491 11509 28503 11543
rect 28445 11503 28503 11509
rect 1104 11450 31280 11472
rect 1104 11398 4182 11450
rect 4234 11398 4246 11450
rect 4298 11398 4310 11450
rect 4362 11398 4374 11450
rect 4426 11398 4438 11450
rect 4490 11398 4502 11450
rect 4554 11398 10182 11450
rect 10234 11398 10246 11450
rect 10298 11398 10310 11450
rect 10362 11398 10374 11450
rect 10426 11398 10438 11450
rect 10490 11398 10502 11450
rect 10554 11398 16182 11450
rect 16234 11398 16246 11450
rect 16298 11398 16310 11450
rect 16362 11398 16374 11450
rect 16426 11398 16438 11450
rect 16490 11398 16502 11450
rect 16554 11398 22182 11450
rect 22234 11398 22246 11450
rect 22298 11398 22310 11450
rect 22362 11398 22374 11450
rect 22426 11398 22438 11450
rect 22490 11398 22502 11450
rect 22554 11398 28182 11450
rect 28234 11398 28246 11450
rect 28298 11398 28310 11450
rect 28362 11398 28374 11450
rect 28426 11398 28438 11450
rect 28490 11398 28502 11450
rect 28554 11398 31280 11450
rect 1104 11376 31280 11398
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 4614 11336 4620 11348
rect 4488 11308 4620 11336
rect 4488 11296 4494 11308
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 10686 11336 10692 11348
rect 10367 11308 10692 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11330 11336 11336 11348
rect 11195 11308 11336 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 11440 11308 13921 11336
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 3651 11240 4568 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 4540 11212 4568 11240
rect 9950 11228 9956 11280
rect 10008 11268 10014 11280
rect 11440 11268 11468 11308
rect 13909 11305 13921 11308
rect 13955 11336 13967 11339
rect 14734 11336 14740 11348
rect 13955 11308 14740 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 17310 11296 17316 11348
rect 17368 11296 17374 11348
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18690 11336 18696 11348
rect 18380 11308 18696 11336
rect 18380 11296 18386 11308
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 21450 11296 21456 11348
rect 21508 11336 21514 11348
rect 21821 11339 21879 11345
rect 21821 11336 21833 11339
rect 21508 11308 21833 11336
rect 21508 11296 21514 11308
rect 21821 11305 21833 11308
rect 21867 11305 21879 11339
rect 21821 11299 21879 11305
rect 26418 11296 26424 11348
rect 26476 11336 26482 11348
rect 26786 11336 26792 11348
rect 26476 11308 26792 11336
rect 26476 11296 26482 11308
rect 26786 11296 26792 11308
rect 26844 11296 26850 11348
rect 26878 11296 26884 11348
rect 26936 11296 26942 11348
rect 27249 11339 27307 11345
rect 27249 11305 27261 11339
rect 27295 11336 27307 11339
rect 27614 11336 27620 11348
rect 27295 11308 27620 11336
rect 27295 11305 27307 11308
rect 27249 11299 27307 11305
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 27706 11296 27712 11348
rect 27764 11296 27770 11348
rect 10008 11240 11468 11268
rect 10008 11228 10014 11240
rect 17862 11228 17868 11280
rect 17920 11268 17926 11280
rect 22646 11268 22652 11280
rect 17920 11240 22140 11268
rect 17920 11228 17926 11240
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 2096 11172 2237 11200
rect 2096 11160 2102 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 4522 11160 4528 11212
rect 4580 11160 4586 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 7984 11172 8953 11200
rect 7984 11160 7990 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11200 10655 11203
rect 10870 11200 10876 11212
rect 10643 11172 10876 11200
rect 10643 11169 10655 11172
rect 10597 11163 10655 11169
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11790 11160 11796 11212
rect 11848 11160 11854 11212
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12526 11200 12532 11212
rect 12483 11172 12532 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 19429 11203 19487 11209
rect 19429 11169 19441 11203
rect 19475 11200 19487 11203
rect 20346 11200 20352 11212
rect 19475 11172 20352 11200
rect 19475 11169 19487 11172
rect 19429 11163 19487 11169
rect 20346 11160 20352 11172
rect 20404 11160 20410 11212
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4764 11104 4997 11132
rect 4764 11092 4770 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 8754 11092 8760 11144
rect 8812 11132 8818 11144
rect 9197 11135 9255 11141
rect 9197 11132 9209 11135
rect 8812 11104 9209 11132
rect 8812 11092 8818 11104
rect 9197 11101 9209 11104
rect 9243 11101 9255 11135
rect 9197 11095 9255 11101
rect 9582 11092 9588 11144
rect 9640 11132 9646 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 9640 11104 10793 11132
rect 9640 11092 9646 11104
rect 10781 11101 10793 11104
rect 10827 11132 10839 11135
rect 10827 11104 12020 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 2492 11067 2550 11073
rect 2492 11033 2504 11067
rect 2538 11064 2550 11067
rect 2958 11064 2964 11076
rect 2538 11036 2964 11064
rect 2538 11033 2550 11036
rect 2492 11027 2550 11033
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 3973 11067 4031 11073
rect 3973 11033 3985 11067
rect 4019 11064 4031 11067
rect 4614 11064 4620 11076
rect 4019 11036 4620 11064
rect 4019 11033 4031 11036
rect 3973 11027 4031 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 10689 11067 10747 11073
rect 10689 11033 10701 11067
rect 10735 11064 10747 11067
rect 11241 11067 11299 11073
rect 11241 11064 11253 11067
rect 10735 11036 11253 11064
rect 10735 11033 10747 11036
rect 10689 11027 10747 11033
rect 11241 11033 11253 11036
rect 11287 11033 11299 11067
rect 11241 11027 11299 11033
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 11790 11064 11796 11076
rect 11480 11036 11796 11064
rect 11480 11024 11486 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 11992 11064 12020 11104
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 15102 11132 15108 11144
rect 14323 11104 15108 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16758 11132 16764 11144
rect 15979 11104 16764 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17218 11092 17224 11144
rect 17276 11132 17282 11144
rect 17276 11104 22048 11132
rect 17276 11092 17282 11104
rect 12710 11064 12716 11076
rect 11992 11036 12716 11064
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 13662 11036 14197 11064
rect 14185 11033 14197 11036
rect 14231 11033 14243 11067
rect 14185 11027 14243 11033
rect 16022 11024 16028 11076
rect 16080 11064 16086 11076
rect 16178 11067 16236 11073
rect 16178 11064 16190 11067
rect 16080 11036 16190 11064
rect 16080 11024 16086 11036
rect 16178 11033 16190 11036
rect 16224 11033 16236 11067
rect 16178 11027 16236 11033
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 20165 11067 20223 11073
rect 20165 11064 20177 11067
rect 19392 11036 20177 11064
rect 19392 11024 19398 11036
rect 20165 11033 20177 11036
rect 20211 11064 20223 11067
rect 21542 11064 21548 11076
rect 20211 11036 21548 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 21542 11024 21548 11036
rect 21600 11024 21606 11076
rect 5626 10956 5632 11008
rect 5684 10956 5690 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 12066 10996 12072 11008
rect 11664 10968 12072 10996
rect 11664 10956 11670 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 22020 10996 22048 11104
rect 22112 11064 22140 11240
rect 22388 11240 22652 11268
rect 22388 11200 22416 11240
rect 22646 11228 22652 11240
rect 22704 11228 22710 11280
rect 22296 11172 22416 11200
rect 22465 11203 22523 11209
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 22296 11132 22324 11172
rect 22465 11169 22477 11203
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 22235 11104 22324 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22480 11132 22508 11163
rect 22428 11104 22508 11132
rect 26697 11135 26755 11141
rect 22428 11092 22434 11104
rect 26697 11101 26709 11135
rect 26743 11132 26755 11135
rect 26896 11132 26924 11296
rect 27724 11200 27752 11296
rect 26988 11172 27752 11200
rect 26988 11141 27016 11172
rect 26743 11104 26924 11132
rect 26973 11135 27031 11141
rect 26743 11101 26755 11104
rect 26697 11095 26755 11101
rect 26973 11101 26985 11135
rect 27019 11101 27031 11135
rect 26973 11095 27031 11101
rect 27065 11135 27123 11141
rect 27065 11101 27077 11135
rect 27111 11132 27123 11135
rect 27154 11132 27160 11144
rect 27111 11104 27160 11132
rect 27111 11101 27123 11104
rect 27065 11095 27123 11101
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 27338 11092 27344 11144
rect 27396 11092 27402 11144
rect 22281 11067 22339 11073
rect 22281 11064 22293 11067
rect 22112 11036 22293 11064
rect 22281 11033 22293 11036
rect 22327 11064 22339 11067
rect 22327 11036 22988 11064
rect 22327 11033 22339 11036
rect 22281 11027 22339 11033
rect 22370 10996 22376 11008
rect 22020 10968 22376 10996
rect 22370 10956 22376 10968
rect 22428 10956 22434 11008
rect 22960 10996 22988 11036
rect 25774 11024 25780 11076
rect 25832 11064 25838 11076
rect 26881 11067 26939 11073
rect 26881 11064 26893 11067
rect 25832 11036 26893 11064
rect 25832 11024 25838 11036
rect 26881 11033 26893 11036
rect 26927 11033 26939 11067
rect 26881 11027 26939 11033
rect 27356 10996 27384 11092
rect 22960 10968 27384 10996
rect 1104 10906 31280 10928
rect 1104 10854 4922 10906
rect 4974 10854 4986 10906
rect 5038 10854 5050 10906
rect 5102 10854 5114 10906
rect 5166 10854 5178 10906
rect 5230 10854 5242 10906
rect 5294 10854 10922 10906
rect 10974 10854 10986 10906
rect 11038 10854 11050 10906
rect 11102 10854 11114 10906
rect 11166 10854 11178 10906
rect 11230 10854 11242 10906
rect 11294 10854 16922 10906
rect 16974 10854 16986 10906
rect 17038 10854 17050 10906
rect 17102 10854 17114 10906
rect 17166 10854 17178 10906
rect 17230 10854 17242 10906
rect 17294 10854 22922 10906
rect 22974 10854 22986 10906
rect 23038 10854 23050 10906
rect 23102 10854 23114 10906
rect 23166 10854 23178 10906
rect 23230 10854 23242 10906
rect 23294 10854 28922 10906
rect 28974 10854 28986 10906
rect 29038 10854 29050 10906
rect 29102 10854 29114 10906
rect 29166 10854 29178 10906
rect 29230 10854 29242 10906
rect 29294 10854 31280 10906
rect 1104 10832 31280 10854
rect 2958 10752 2964 10804
rect 3016 10752 3022 10804
rect 4706 10752 4712 10804
rect 4764 10752 4770 10804
rect 4798 10752 4804 10804
rect 4856 10752 4862 10804
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5626 10792 5632 10804
rect 5215 10764 5632 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 9861 10795 9919 10801
rect 9861 10792 9873 10795
rect 9732 10764 9873 10792
rect 9732 10752 9738 10764
rect 9861 10761 9873 10764
rect 9907 10761 9919 10795
rect 9861 10755 9919 10761
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 25774 10792 25780 10804
rect 24811 10764 25780 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 3596 10727 3654 10733
rect 3596 10693 3608 10727
rect 3642 10724 3654 10727
rect 3786 10724 3792 10736
rect 3642 10696 3792 10724
rect 3642 10693 3654 10696
rect 3596 10687 3654 10693
rect 3786 10684 3792 10696
rect 3844 10684 3850 10736
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 5261 10727 5319 10733
rect 5261 10724 5273 10727
rect 4120 10696 5273 10724
rect 4120 10684 4126 10696
rect 5261 10693 5273 10696
rect 5307 10724 5319 10727
rect 5307 10696 6960 10724
rect 5307 10693 5319 10696
rect 5261 10687 5319 10693
rect 3142 10616 3148 10668
rect 3200 10616 3206 10668
rect 3970 10656 3976 10668
rect 3252 10628 3976 10656
rect 3252 10600 3280 10628
rect 3970 10616 3976 10628
rect 4028 10656 4034 10668
rect 4028 10628 5396 10656
rect 4028 10616 4034 10628
rect 3234 10548 3240 10600
rect 3292 10548 3298 10600
rect 3326 10548 3332 10600
rect 3384 10548 3390 10600
rect 5368 10597 5396 10628
rect 6932 10600 6960 10696
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10686 10656 10692 10668
rect 10551 10628 10692 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 23900 10628 24409 10656
rect 23900 10616 23906 10628
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10557 5411 10591
rect 5353 10551 5411 10557
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 24486 10548 24492 10600
rect 24544 10548 24550 10600
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 4798 10520 4804 10532
rect 4580 10492 4804 10520
rect 4580 10480 4586 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4890 10452 4896 10464
rect 4488 10424 4896 10452
rect 4488 10412 4494 10424
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 24397 10455 24455 10461
rect 24397 10452 24409 10455
rect 21968 10424 24409 10452
rect 21968 10412 21974 10424
rect 24397 10421 24409 10424
rect 24443 10421 24455 10455
rect 24397 10415 24455 10421
rect 1104 10362 31280 10384
rect 1104 10310 4182 10362
rect 4234 10310 4246 10362
rect 4298 10310 4310 10362
rect 4362 10310 4374 10362
rect 4426 10310 4438 10362
rect 4490 10310 4502 10362
rect 4554 10310 10182 10362
rect 10234 10310 10246 10362
rect 10298 10310 10310 10362
rect 10362 10310 10374 10362
rect 10426 10310 10438 10362
rect 10490 10310 10502 10362
rect 10554 10310 16182 10362
rect 16234 10310 16246 10362
rect 16298 10310 16310 10362
rect 16362 10310 16374 10362
rect 16426 10310 16438 10362
rect 16490 10310 16502 10362
rect 16554 10310 22182 10362
rect 22234 10310 22246 10362
rect 22298 10310 22310 10362
rect 22362 10310 22374 10362
rect 22426 10310 22438 10362
rect 22490 10310 22502 10362
rect 22554 10310 28182 10362
rect 28234 10310 28246 10362
rect 28298 10310 28310 10362
rect 28362 10310 28374 10362
rect 28426 10310 28438 10362
rect 28490 10310 28502 10362
rect 28554 10310 31280 10362
rect 1104 10288 31280 10310
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3200 10220 3801 10248
rect 3200 10208 3206 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 5442 10248 5448 10260
rect 4120 10220 4200 10248
rect 4120 10208 4126 10220
rect 4172 10112 4200 10220
rect 4356 10220 5448 10248
rect 4356 10124 4384 10220
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 23566 10208 23572 10260
rect 23624 10208 23630 10260
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 4172 10084 4261 10112
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4249 10075 4307 10081
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 4724 10084 5120 10112
rect 4724 10056 4752 10084
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4614 10044 4620 10056
rect 4203 10016 4620 10044
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5092 10053 5120 10084
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19978 10112 19984 10124
rect 19484 10084 19984 10112
rect 19484 10072 19490 10084
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 22554 10072 22560 10124
rect 22612 10112 22618 10124
rect 22612 10084 23336 10112
rect 22612 10072 22618 10084
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4948 10016 4997 10044
rect 4948 10004 4954 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5350 10044 5356 10056
rect 5215 10016 5356 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 7742 10004 7748 10056
rect 7800 10004 7806 10056
rect 9950 10004 9956 10056
rect 10008 10044 10014 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 10008 10016 10425 10044
rect 10008 10004 10014 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 20806 10004 20812 10056
rect 20864 10004 20870 10056
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 23308 10053 23336 10084
rect 22925 10047 22983 10053
rect 22925 10044 22937 10047
rect 22428 10016 22937 10044
rect 22428 10004 22434 10016
rect 22925 10013 22937 10016
rect 22971 10013 22983 10047
rect 22925 10007 22983 10013
rect 23293 10047 23351 10053
rect 23293 10013 23305 10047
rect 23339 10044 23351 10047
rect 23584 10044 23612 10208
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25961 10115 26019 10121
rect 25961 10112 25973 10115
rect 25004 10084 25973 10112
rect 25004 10072 25010 10084
rect 25961 10081 25973 10084
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 23339 10016 23612 10044
rect 23339 10013 23351 10016
rect 23293 10007 23351 10013
rect 25038 10004 25044 10056
rect 25096 10044 25102 10056
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 25096 10016 25237 10044
rect 25096 10004 25102 10016
rect 25225 10013 25237 10016
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 4908 9908 4936 10004
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 20257 9979 20315 9985
rect 20257 9976 20269 9979
rect 19843 9948 20269 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 20257 9945 20269 9948
rect 20303 9945 20315 9979
rect 20257 9939 20315 9945
rect 22738 9936 22744 9988
rect 22796 9976 22802 9988
rect 23109 9979 23167 9985
rect 23109 9976 23121 9979
rect 22796 9948 23121 9976
rect 22796 9936 22802 9948
rect 23109 9945 23121 9948
rect 23155 9945 23167 9979
rect 23109 9939 23167 9945
rect 23201 9979 23259 9985
rect 23201 9945 23213 9979
rect 23247 9976 23259 9979
rect 23566 9976 23572 9988
rect 23247 9948 23572 9976
rect 23247 9945 23259 9948
rect 23201 9939 23259 9945
rect 23566 9936 23572 9948
rect 23624 9936 23630 9988
rect 4856 9880 4936 9908
rect 5353 9911 5411 9917
rect 4856 9868 4862 9880
rect 5353 9877 5365 9911
rect 5399 9908 5411 9911
rect 6362 9908 6368 9920
rect 5399 9880 6368 9908
rect 5399 9877 5411 9880
rect 5353 9871 5411 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7190 9868 7196 9920
rect 7248 9868 7254 9920
rect 9858 9868 9864 9920
rect 9916 9868 9922 9920
rect 17402 9868 17408 9920
rect 17460 9868 17466 9920
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19429 9911 19487 9917
rect 19429 9908 19441 9911
rect 19392 9880 19441 9908
rect 19392 9868 19398 9880
rect 19429 9877 19441 9880
rect 19475 9877 19487 9911
rect 19429 9871 19487 9877
rect 19610 9868 19616 9920
rect 19668 9908 19674 9920
rect 19889 9911 19947 9917
rect 19889 9908 19901 9911
rect 19668 9880 19901 9908
rect 19668 9868 19674 9880
rect 19889 9877 19901 9880
rect 19935 9877 19947 9911
rect 19889 9871 19947 9877
rect 23474 9868 23480 9920
rect 23532 9868 23538 9920
rect 24210 9868 24216 9920
rect 24268 9908 24274 9920
rect 24578 9908 24584 9920
rect 24268 9880 24584 9908
rect 24268 9868 24274 9880
rect 24578 9868 24584 9880
rect 24636 9868 24642 9920
rect 24673 9911 24731 9917
rect 24673 9877 24685 9911
rect 24719 9908 24731 9911
rect 24854 9908 24860 9920
rect 24719 9880 24860 9908
rect 24719 9877 24731 9880
rect 24673 9871 24731 9877
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 25406 9868 25412 9920
rect 25464 9868 25470 9920
rect 1104 9818 31280 9840
rect 1104 9766 4922 9818
rect 4974 9766 4986 9818
rect 5038 9766 5050 9818
rect 5102 9766 5114 9818
rect 5166 9766 5178 9818
rect 5230 9766 5242 9818
rect 5294 9766 10922 9818
rect 10974 9766 10986 9818
rect 11038 9766 11050 9818
rect 11102 9766 11114 9818
rect 11166 9766 11178 9818
rect 11230 9766 11242 9818
rect 11294 9766 16922 9818
rect 16974 9766 16986 9818
rect 17038 9766 17050 9818
rect 17102 9766 17114 9818
rect 17166 9766 17178 9818
rect 17230 9766 17242 9818
rect 17294 9766 22922 9818
rect 22974 9766 22986 9818
rect 23038 9766 23050 9818
rect 23102 9766 23114 9818
rect 23166 9766 23178 9818
rect 23230 9766 23242 9818
rect 23294 9766 28922 9818
rect 28974 9766 28986 9818
rect 29038 9766 29050 9818
rect 29102 9766 29114 9818
rect 29166 9766 29178 9818
rect 29230 9766 29242 9818
rect 29294 9766 31280 9818
rect 1104 9744 31280 9766
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9704 6975 9707
rect 7190 9704 7196 9716
rect 6963 9676 7196 9704
rect 6963 9673 6975 9676
rect 6917 9667 6975 9673
rect 7190 9664 7196 9676
rect 7248 9664 7254 9716
rect 9677 9707 9735 9713
rect 9677 9673 9689 9707
rect 9723 9704 9735 9707
rect 9858 9704 9864 9716
rect 9723 9676 9864 9704
rect 9723 9673 9735 9676
rect 9677 9667 9735 9673
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 17129 9707 17187 9713
rect 17129 9673 17141 9707
rect 17175 9704 17187 9707
rect 17402 9704 17408 9716
rect 17175 9676 17408 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17402 9664 17408 9676
rect 17460 9664 17466 9716
rect 21361 9707 21419 9713
rect 21361 9673 21373 9707
rect 21407 9704 21419 9707
rect 21407 9676 21441 9704
rect 21407 9673 21419 9676
rect 21361 9667 21419 9673
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 7098 9636 7104 9648
rect 7055 9608 7104 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 7098 9596 7104 9608
rect 7156 9596 7162 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7653 9639 7711 9645
rect 7653 9636 7665 9639
rect 7340 9608 7665 9636
rect 7340 9596 7346 9608
rect 7653 9605 7665 9608
rect 7699 9636 7711 9639
rect 8294 9636 8300 9648
rect 7699 9608 8300 9636
rect 7699 9605 7711 9608
rect 7653 9599 7711 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9217 9639 9275 9645
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 10413 9639 10471 9645
rect 10413 9636 10425 9639
rect 9263 9608 10425 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 10413 9605 10425 9608
rect 10459 9636 10471 9639
rect 15378 9636 15384 9648
rect 10459 9608 15384 9636
rect 10459 9605 10471 9608
rect 10413 9599 10471 9605
rect 15378 9596 15384 9608
rect 15436 9636 15442 9648
rect 18322 9636 18328 9648
rect 15436 9608 18328 9636
rect 15436 9596 15442 9608
rect 18322 9596 18328 9608
rect 18380 9636 18386 9648
rect 19242 9636 19248 9648
rect 18380 9608 19248 9636
rect 18380 9596 18386 9608
rect 19242 9596 19248 9608
rect 19300 9596 19306 9648
rect 21376 9636 21404 9667
rect 21910 9664 21916 9716
rect 21968 9664 21974 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 23382 9704 23388 9716
rect 22428 9676 23388 9704
rect 22428 9664 22434 9676
rect 23382 9664 23388 9676
rect 23440 9664 23446 9716
rect 23750 9704 23756 9716
rect 23584 9676 23756 9704
rect 21928 9636 21956 9664
rect 22465 9639 22523 9645
rect 22465 9636 22477 9639
rect 21376 9608 21956 9636
rect 22066 9608 22477 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2961 9571 3019 9577
rect 2547 9540 2636 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2608 9441 2636 9540
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3007 9540 3433 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 5718 9568 5724 9580
rect 3844 9540 5724 9568
rect 3844 9528 3850 9540
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 7558 9577 7564 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 6420 9540 7389 9568
rect 6420 9528 6426 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7525 9571 7564 9577
rect 7525 9537 7537 9571
rect 7525 9531 7564 9537
rect 7558 9528 7564 9531
rect 7616 9528 7622 9580
rect 7742 9528 7748 9580
rect 7800 9528 7806 9580
rect 7834 9528 7840 9580
rect 7892 9577 7898 9580
rect 7892 9568 7900 9577
rect 8478 9568 8484 9580
rect 7892 9540 8484 9568
rect 7892 9531 7900 9540
rect 7892 9528 7898 9531
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11112 9540 11253 9568
rect 11112 9528 11118 9540
rect 11241 9537 11253 9540
rect 11287 9568 11299 9571
rect 12158 9568 12164 9580
rect 11287 9540 12164 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12250 9528 12256 9580
rect 12308 9528 12314 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9568 15991 9571
rect 18049 9571 18107 9577
rect 15979 9540 16804 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9500 4123 9503
rect 4111 9472 4752 9500
rect 4111 9469 4123 9472
rect 4065 9463 4123 9469
rect 2593 9435 2651 9441
rect 2593 9401 2605 9435
rect 2639 9401 2651 9435
rect 2593 9395 2651 9401
rect 2314 9324 2320 9376
rect 2372 9324 2378 9376
rect 3068 9364 3096 9463
rect 3160 9432 3188 9463
rect 4338 9432 4344 9444
rect 3160 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 4724 9376 4752 9472
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7101 9503 7159 9509
rect 7101 9500 7113 9503
rect 6880 9472 7113 9500
rect 6880 9460 6886 9472
rect 7101 9469 7113 9472
rect 7147 9469 7159 9503
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 7101 9463 7159 9469
rect 7300 9472 8401 9500
rect 6012 9404 6776 9432
rect 6012 9376 6040 9404
rect 3786 9364 3792 9376
rect 3068 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 5994 9324 6000 9376
rect 6052 9324 6058 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 6748 9364 6776 9404
rect 7300 9364 7328 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 9769 9503 9827 9509
rect 9769 9469 9781 9503
rect 9815 9500 9827 9503
rect 9858 9500 9864 9512
rect 9815 9472 9864 9500
rect 9815 9469 9827 9472
rect 9769 9463 9827 9469
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10042 9500 10048 9512
rect 9999 9472 10048 9500
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11020 9472 12081 9500
rect 11020 9460 11026 9472
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 12342 9460 12348 9512
rect 12400 9460 12406 9512
rect 16776 9441 16804 9540
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18095 9540 18521 9568
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19501 9571 19559 9577
rect 19501 9568 19513 9571
rect 19208 9540 19513 9568
rect 19208 9528 19214 9540
rect 19501 9537 19513 9540
rect 19547 9537 19559 9571
rect 19501 9531 19559 9537
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 19944 9540 20729 9568
rect 19944 9528 19950 9540
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20806 9528 20812 9580
rect 20864 9568 20870 9580
rect 20864 9540 20909 9568
rect 20864 9528 20870 9540
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 21082 9528 21088 9580
rect 21140 9528 21146 9580
rect 21174 9528 21180 9580
rect 21232 9577 21238 9580
rect 21232 9531 21240 9577
rect 21232 9528 21238 9531
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 16761 9435 16819 9441
rect 9232 9404 12296 9432
rect 6748 9336 7328 9364
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 9232 9364 9260 9404
rect 8067 9336 9260 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 9306 9324 9312 9376
rect 9364 9324 9370 9376
rect 11514 9324 11520 9376
rect 11572 9324 11578 9376
rect 12268 9373 12296 9404
rect 16761 9401 16773 9435
rect 16807 9401 16819 9435
rect 17236 9432 17264 9463
rect 17310 9460 17316 9512
rect 17368 9460 17374 9512
rect 18141 9503 18199 9509
rect 18141 9469 18153 9503
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 18156 9432 18184 9463
rect 17236 9404 18184 9432
rect 16761 9395 16819 9401
rect 12253 9367 12311 9373
rect 12253 9333 12265 9367
rect 12299 9333 12311 9367
rect 12253 9327 12311 9333
rect 12618 9324 12624 9376
rect 12676 9324 12682 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 16080 9336 16129 9364
rect 16080 9324 16086 9336
rect 16117 9333 16129 9336
rect 16163 9333 16175 9367
rect 16117 9327 16175 9333
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 16632 9336 17693 9364
rect 16632 9324 16638 9336
rect 17681 9333 17693 9336
rect 17727 9333 17739 9367
rect 18156 9364 18184 9404
rect 18230 9392 18236 9444
rect 18288 9432 18294 9444
rect 18340 9432 18368 9463
rect 19058 9460 19064 9512
rect 19116 9460 19122 9512
rect 19242 9460 19248 9512
rect 19300 9460 19306 9512
rect 18288 9404 18368 9432
rect 20625 9435 20683 9441
rect 18288 9392 18294 9404
rect 20625 9401 20637 9435
rect 20671 9432 20683 9435
rect 20824 9432 20852 9528
rect 20898 9460 20904 9512
rect 20956 9500 20962 9512
rect 21197 9500 21225 9528
rect 20956 9472 21225 9500
rect 20956 9460 20962 9472
rect 22066 9432 22094 9608
rect 22465 9605 22477 9608
rect 22511 9636 22523 9639
rect 23584 9636 23612 9676
rect 23750 9664 23756 9676
rect 23808 9704 23814 9716
rect 24397 9707 24455 9713
rect 23808 9676 24348 9704
rect 23808 9664 23814 9676
rect 22511 9608 23612 9636
rect 22511 9605 22523 9608
rect 22465 9599 22523 9605
rect 23658 9596 23664 9648
rect 23716 9636 23722 9648
rect 24121 9639 24179 9645
rect 23716 9608 24072 9636
rect 23716 9596 23722 9608
rect 24044 9580 24072 9608
rect 24121 9605 24133 9639
rect 24167 9605 24179 9639
rect 24320 9636 24348 9676
rect 24397 9673 24409 9707
rect 24443 9704 24455 9707
rect 24486 9704 24492 9716
rect 24443 9676 24492 9704
rect 24443 9673 24455 9676
rect 24397 9667 24455 9673
rect 24486 9664 24492 9676
rect 24544 9664 24550 9716
rect 24765 9707 24823 9713
rect 24765 9673 24777 9707
rect 24811 9704 24823 9707
rect 24854 9704 24860 9716
rect 24811 9676 24860 9704
rect 24811 9673 24823 9676
rect 24765 9667 24823 9673
rect 24854 9664 24860 9676
rect 24912 9664 24918 9716
rect 24964 9676 25176 9704
rect 24964 9636 24992 9676
rect 24320 9608 24992 9636
rect 25148 9636 25176 9676
rect 25406 9664 25412 9716
rect 25464 9704 25470 9716
rect 25593 9707 25651 9713
rect 25593 9704 25605 9707
rect 25464 9676 25605 9704
rect 25464 9664 25470 9676
rect 25593 9673 25605 9676
rect 25639 9673 25651 9707
rect 25593 9667 25651 9673
rect 25148 9608 26188 9636
rect 24121 9599 24179 9605
rect 22373 9571 22431 9577
rect 22373 9537 22385 9571
rect 22419 9568 22431 9571
rect 22833 9571 22891 9577
rect 22833 9568 22845 9571
rect 22419 9540 22845 9568
rect 22419 9537 22431 9540
rect 22373 9531 22431 9537
rect 22833 9537 22845 9540
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 23382 9528 23388 9580
rect 23440 9528 23446 9580
rect 23474 9528 23480 9580
rect 23532 9568 23538 9580
rect 23753 9571 23811 9577
rect 23753 9568 23765 9571
rect 23532 9540 23765 9568
rect 23532 9528 23538 9540
rect 23753 9537 23765 9540
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 23901 9571 23959 9577
rect 23901 9537 23913 9571
rect 23947 9568 23959 9571
rect 23947 9537 23980 9568
rect 23901 9531 23980 9537
rect 22646 9460 22652 9512
rect 22704 9460 22710 9512
rect 20671 9404 20852 9432
rect 20916 9404 22094 9432
rect 20671 9401 20683 9404
rect 20625 9395 20683 9401
rect 20916 9364 20944 9404
rect 18156 9336 20944 9364
rect 17681 9327 17739 9333
rect 22002 9324 22008 9376
rect 22060 9324 22066 9376
rect 23952 9364 23980 9531
rect 24026 9528 24032 9580
rect 24084 9528 24090 9580
rect 24136 9444 24164 9599
rect 24218 9571 24276 9577
rect 24218 9537 24230 9571
rect 24264 9537 24276 9571
rect 24218 9531 24276 9537
rect 24118 9392 24124 9444
rect 24176 9392 24182 9444
rect 24228 9432 24256 9531
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 26160 9577 26188 9608
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24820 9540 24869 9568
rect 24820 9528 24826 9540
rect 24857 9537 24869 9540
rect 24903 9568 24915 9571
rect 25685 9571 25743 9577
rect 25685 9568 25697 9571
rect 24903 9540 25697 9568
rect 24903 9537 24915 9540
rect 24857 9531 24915 9537
rect 25685 9537 25697 9540
rect 25731 9568 25743 9571
rect 26145 9571 26203 9577
rect 25731 9540 26004 9568
rect 25731 9537 25743 9540
rect 25685 9531 25743 9537
rect 24394 9460 24400 9512
rect 24452 9500 24458 9512
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 24452 9472 24593 9500
rect 24452 9460 24458 9472
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 25406 9460 25412 9512
rect 25464 9500 25470 9512
rect 25866 9500 25872 9512
rect 25464 9472 25872 9500
rect 25464 9460 25470 9472
rect 25866 9460 25872 9472
rect 25924 9460 25930 9512
rect 25976 9500 26004 9540
rect 26145 9537 26157 9571
rect 26191 9568 26203 9571
rect 30742 9568 30748 9580
rect 26191 9540 30748 9568
rect 26191 9537 26203 9540
rect 26145 9531 26203 9537
rect 30742 9528 30748 9540
rect 30800 9528 30806 9580
rect 26418 9500 26424 9512
rect 25976 9472 26424 9500
rect 26418 9460 26424 9472
rect 26476 9460 26482 9512
rect 24302 9432 24308 9444
rect 24228 9404 24308 9432
rect 24302 9392 24308 9404
rect 24360 9432 24366 9444
rect 24854 9432 24860 9444
rect 24360 9404 24860 9432
rect 24360 9392 24366 9404
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 24946 9392 24952 9444
rect 25004 9392 25010 9444
rect 26329 9435 26387 9441
rect 26329 9401 26341 9435
rect 26375 9432 26387 9435
rect 26436 9432 26464 9460
rect 26375 9404 26464 9432
rect 26375 9401 26387 9404
rect 26329 9395 26387 9401
rect 24964 9364 24992 9392
rect 23952 9336 24992 9364
rect 25225 9367 25283 9373
rect 25225 9333 25237 9367
rect 25271 9364 25283 9367
rect 25590 9364 25596 9376
rect 25271 9336 25596 9364
rect 25271 9333 25283 9336
rect 25225 9327 25283 9333
rect 25590 9324 25596 9336
rect 25648 9324 25654 9376
rect 26050 9324 26056 9376
rect 26108 9324 26114 9376
rect 1104 9274 31280 9296
rect 1104 9222 4182 9274
rect 4234 9222 4246 9274
rect 4298 9222 4310 9274
rect 4362 9222 4374 9274
rect 4426 9222 4438 9274
rect 4490 9222 4502 9274
rect 4554 9222 10182 9274
rect 10234 9222 10246 9274
rect 10298 9222 10310 9274
rect 10362 9222 10374 9274
rect 10426 9222 10438 9274
rect 10490 9222 10502 9274
rect 10554 9222 16182 9274
rect 16234 9222 16246 9274
rect 16298 9222 16310 9274
rect 16362 9222 16374 9274
rect 16426 9222 16438 9274
rect 16490 9222 16502 9274
rect 16554 9222 22182 9274
rect 22234 9222 22246 9274
rect 22298 9222 22310 9274
rect 22362 9222 22374 9274
rect 22426 9222 22438 9274
rect 22490 9222 22502 9274
rect 22554 9222 28182 9274
rect 28234 9222 28246 9274
rect 28298 9222 28310 9274
rect 28362 9222 28374 9274
rect 28426 9222 28438 9274
rect 28490 9222 28502 9274
rect 28554 9222 31280 9274
rect 1104 9200 31280 9222
rect 5828 9132 6040 9160
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 4706 9092 4712 9104
rect 3375 9064 4712 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 5828 9024 5856 9132
rect 5905 9095 5963 9101
rect 5905 9061 5917 9095
rect 5951 9061 5963 9095
rect 5905 9055 5963 9061
rect 3344 8996 5856 9024
rect 3344 8968 3372 8996
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2774 8956 2780 8968
rect 1995 8928 2780 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2774 8916 2780 8928
rect 2832 8956 2838 8968
rect 3326 8956 3332 8968
rect 2832 8928 3332 8956
rect 2832 8916 2838 8928
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 5920 8956 5948 9055
rect 6012 9036 6040 9132
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6638 9160 6644 9172
rect 6236 9132 6644 9160
rect 6236 9120 6242 9132
rect 6638 9120 6644 9132
rect 6696 9160 6702 9172
rect 7377 9163 7435 9169
rect 6696 9132 7052 9160
rect 6696 9120 6702 9132
rect 5994 8984 6000 9036
rect 6052 8984 6058 9036
rect 7024 9024 7052 9132
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7742 9160 7748 9172
rect 7423 9132 7748 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 9306 9120 9312 9172
rect 9364 9120 9370 9172
rect 12253 9163 12311 9169
rect 10520 9132 12204 9160
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7024 8996 8033 9024
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 9324 9024 9352 9120
rect 10520 9036 10548 9132
rect 10873 9095 10931 9101
rect 10873 9061 10885 9095
rect 10919 9092 10931 9095
rect 10962 9092 10968 9104
rect 10919 9064 10968 9092
rect 10919 9061 10931 9064
rect 10873 9055 10931 9061
rect 10962 9052 10968 9064
rect 11020 9092 11026 9104
rect 12176 9092 12204 9132
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12342 9160 12348 9172
rect 12299 9132 12348 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 19061 9163 19119 9169
rect 19061 9129 19073 9163
rect 19107 9160 19119 9163
rect 19150 9160 19156 9172
rect 19107 9132 19156 9160
rect 19107 9129 19119 9132
rect 19061 9123 19119 9129
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19242 9120 19248 9172
rect 19300 9120 19306 9172
rect 19610 9120 19616 9172
rect 19668 9160 19674 9172
rect 20625 9163 20683 9169
rect 19668 9132 20576 9160
rect 19668 9120 19674 9132
rect 11020 9064 11192 9092
rect 12176 9064 12756 9092
rect 11020 9052 11026 9064
rect 8021 8987 8079 8993
rect 9140 8996 9352 9024
rect 6253 8959 6311 8965
rect 6253 8956 6265 8959
rect 5767 8928 5856 8956
rect 5920 8928 6265 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 2216 8891 2274 8897
rect 2216 8857 2228 8891
rect 2262 8888 2274 8891
rect 2314 8888 2320 8900
rect 2262 8860 2320 8888
rect 2262 8857 2274 8860
rect 2216 8851 2274 8857
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 4632 8832 4660 8919
rect 5460 8888 5488 8919
rect 5828 8888 5856 8928
rect 6253 8925 6265 8928
rect 6299 8925 6311 8959
rect 6253 8919 6311 8925
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7926 8956 7932 8968
rect 7156 8928 7932 8956
rect 7156 8916 7162 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 9140 8965 9168 8996
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 11054 9024 11060 9036
rect 10612 8996 11060 9024
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 9324 8928 9505 8956
rect 6564 8888 6592 8916
rect 5460 8860 5764 8888
rect 5828 8860 6592 8888
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 4614 8780 4620 8832
rect 4672 8780 4678 8832
rect 5626 8780 5632 8832
rect 5684 8780 5690 8832
rect 5736 8820 5764 8860
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 9324 8888 9352 8928
rect 9493 8925 9505 8928
rect 9539 8956 9551 8959
rect 10612 8956 10640 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11164 9024 11192 9064
rect 12526 9024 12532 9036
rect 11164 8996 11284 9024
rect 9539 8928 10640 8956
rect 10965 8959 11023 8965
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 9738 8891 9796 8897
rect 9738 8888 9750 8891
rect 8720 8860 9352 8888
rect 9416 8860 9750 8888
rect 8720 8848 8726 8860
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 5736 8792 7481 8820
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 7834 8780 7840 8832
rect 7892 8780 7898 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9416 8829 9444 8860
rect 9738 8857 9750 8860
rect 9784 8857 9796 8891
rect 9738 8851 9796 8857
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10980 8888 11008 8919
rect 11146 8916 11152 8968
rect 11204 8916 11210 8968
rect 10008 8860 11008 8888
rect 10008 8848 10014 8860
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8904 8792 8953 8820
rect 8904 8780 8910 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9401 8823 9459 8829
rect 9401 8789 9413 8823
rect 9447 8789 9459 8823
rect 11164 8820 11192 8916
rect 11256 8897 11284 8996
rect 11992 8996 12532 9024
rect 11330 8916 11336 8968
rect 11388 8916 11394 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11532 8928 11621 8956
rect 11241 8891 11299 8897
rect 11241 8857 11253 8891
rect 11287 8857 11299 8891
rect 11241 8851 11299 8857
rect 11422 8820 11428 8832
rect 11164 8792 11428 8820
rect 9401 8783 9459 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 11532 8829 11560 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11757 8959 11815 8965
rect 11757 8925 11769 8959
rect 11803 8956 11815 8959
rect 11992 8956 12020 8996
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 11803 8928 12020 8956
rect 11803 8925 11815 8928
rect 11757 8919 11815 8925
rect 12066 8916 12072 8968
rect 12124 8965 12130 8968
rect 12728 8965 12756 9064
rect 12894 8984 12900 9036
rect 12952 8984 12958 9036
rect 13814 9024 13820 9036
rect 13280 8996 13820 9024
rect 12124 8956 12132 8965
rect 12713 8959 12771 8965
rect 12124 8928 12169 8956
rect 12124 8919 12132 8928
rect 12713 8925 12725 8959
rect 12759 8956 12771 8959
rect 13280 8956 13308 8996
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 19260 9033 19288 9120
rect 20548 9092 20576 9132
rect 20625 9129 20637 9163
rect 20671 9160 20683 9163
rect 21082 9160 21088 9172
rect 20671 9132 21088 9160
rect 20671 9129 20683 9132
rect 20625 9123 20683 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 23109 9163 23167 9169
rect 21192 9132 23060 9160
rect 21192 9092 21220 9132
rect 20548 9064 21220 9092
rect 23032 9092 23060 9132
rect 23109 9129 23121 9163
rect 23155 9160 23167 9163
rect 23382 9160 23388 9172
rect 23155 9132 23388 9160
rect 23155 9129 23167 9132
rect 23109 9123 23167 9129
rect 23382 9120 23388 9132
rect 23440 9120 23446 9172
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24397 9163 24455 9169
rect 24397 9160 24409 9163
rect 24176 9132 24409 9160
rect 24176 9120 24182 9132
rect 24397 9129 24409 9132
rect 24443 9160 24455 9163
rect 25038 9160 25044 9172
rect 24443 9132 25044 9160
rect 24443 9129 24455 9132
rect 24397 9123 24455 9129
rect 25038 9120 25044 9132
rect 25096 9120 25102 9172
rect 25590 9120 25596 9172
rect 25648 9160 25654 9172
rect 25648 9132 26004 9160
rect 25648 9120 25654 9132
rect 23937 9095 23995 9101
rect 23032 9064 23612 9092
rect 19245 9027 19303 9033
rect 19245 8993 19257 9027
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 23293 9027 23351 9033
rect 23293 8993 23305 9027
rect 23339 8993 23351 9027
rect 23293 8987 23351 8993
rect 12759 8928 13308 8956
rect 13725 8959 13783 8965
rect 12759 8925 12771 8928
rect 12713 8919 12771 8925
rect 13725 8925 13737 8959
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 12124 8916 12130 8919
rect 11885 8891 11943 8897
rect 11885 8888 11897 8891
rect 11716 8860 11897 8888
rect 11716 8832 11744 8860
rect 11885 8857 11897 8860
rect 11931 8857 11943 8891
rect 11885 8851 11943 8857
rect 11977 8891 12035 8897
rect 11977 8857 11989 8891
rect 12023 8888 12035 8891
rect 13354 8888 13360 8900
rect 12023 8860 13360 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 13354 8848 13360 8860
rect 13412 8888 13418 8900
rect 13740 8888 13768 8919
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16025 8959 16083 8965
rect 16025 8956 16037 8959
rect 15988 8928 16037 8956
rect 15988 8916 15994 8928
rect 16025 8925 16037 8928
rect 16071 8925 16083 8959
rect 16025 8919 16083 8925
rect 16209 8959 16267 8965
rect 16209 8925 16221 8959
rect 16255 8956 16267 8959
rect 17954 8956 17960 8968
rect 16255 8928 17960 8956
rect 16255 8925 16267 8928
rect 16209 8919 16267 8925
rect 13412 8860 13768 8888
rect 13412 8848 13418 8860
rect 14826 8848 14832 8900
rect 14884 8888 14890 8900
rect 16224 8888 16252 8919
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 18380 8928 18797 8956
rect 18380 8916 18386 8928
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 19150 8956 19156 8968
rect 18923 8928 19156 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 16454 8891 16512 8897
rect 16454 8888 16466 8891
rect 14884 8860 16252 8888
rect 16316 8860 16466 8888
rect 14884 8848 14890 8860
rect 11517 8823 11575 8829
rect 11517 8789 11529 8823
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 11698 8780 11704 8832
rect 11756 8780 11762 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 11848 8792 12357 8820
rect 11848 8780 11854 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 12805 8823 12863 8829
rect 12805 8789 12817 8823
rect 12851 8820 12863 8823
rect 13173 8823 13231 8829
rect 13173 8820 13185 8823
rect 12851 8792 13185 8820
rect 12851 8789 12863 8792
rect 12805 8783 12863 8789
rect 13173 8789 13185 8792
rect 13219 8789 13231 8823
rect 13173 8783 13231 8789
rect 15470 8780 15476 8832
rect 15528 8780 15534 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16316 8820 16344 8860
rect 16454 8857 16466 8860
rect 16500 8857 16512 8891
rect 16454 8851 16512 8857
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17494 8888 17500 8900
rect 16724 8860 17500 8888
rect 16724 8848 16730 8860
rect 17494 8848 17500 8860
rect 17552 8888 17558 8900
rect 18230 8888 18236 8900
rect 17552 8860 18236 8888
rect 17552 8848 17558 8860
rect 18230 8848 18236 8860
rect 18288 8848 18294 8900
rect 18800 8888 18828 8919
rect 19150 8916 19156 8928
rect 19208 8916 19214 8968
rect 19260 8956 19288 8987
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 19260 8928 20821 8956
rect 20809 8925 20821 8928
rect 20855 8956 20867 8959
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 20855 8928 21741 8956
rect 20855 8925 20867 8928
rect 20809 8919 20867 8925
rect 21729 8925 21741 8928
rect 21775 8956 21787 8959
rect 23308 8956 23336 8987
rect 23382 8956 23388 8968
rect 21775 8928 22094 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 19512 8891 19570 8897
rect 18800 8860 19288 8888
rect 16080 8792 16344 8820
rect 17589 8823 17647 8829
rect 16080 8780 16086 8792
rect 17589 8789 17601 8823
rect 17635 8820 17647 8823
rect 18046 8820 18052 8832
rect 17635 8792 18052 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 18046 8780 18052 8792
rect 18104 8820 18110 8832
rect 18782 8820 18788 8832
rect 18104 8792 18788 8820
rect 18104 8780 18110 8792
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19260 8820 19288 8860
rect 19512 8857 19524 8891
rect 19558 8888 19570 8891
rect 20162 8888 20168 8900
rect 19558 8860 20168 8888
rect 19558 8857 19570 8860
rect 19512 8851 19570 8857
rect 20162 8848 20168 8860
rect 20220 8848 20226 8900
rect 21637 8891 21695 8897
rect 21637 8888 21649 8891
rect 20272 8860 21649 8888
rect 20272 8820 20300 8860
rect 21637 8857 21649 8860
rect 21683 8857 21695 8891
rect 21637 8851 21695 8857
rect 21818 8848 21824 8900
rect 21876 8888 21882 8900
rect 21974 8891 22032 8897
rect 21974 8888 21986 8891
rect 21876 8860 21986 8888
rect 21876 8848 21882 8860
rect 21974 8857 21986 8860
rect 22020 8857 22032 8891
rect 21974 8851 22032 8857
rect 19260 8792 20300 8820
rect 22066 8832 22094 8928
rect 22204 8928 23388 8956
rect 22204 8900 22232 8928
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 22186 8848 22192 8900
rect 22244 8848 22250 8900
rect 23584 8897 23612 9064
rect 23937 9061 23949 9095
rect 23983 9061 23995 9095
rect 23937 9055 23995 9061
rect 23952 8956 23980 9055
rect 24026 9052 24032 9104
rect 24084 9092 24090 9104
rect 24578 9092 24584 9104
rect 24084 9064 24584 9092
rect 24084 9052 24090 9064
rect 24578 9052 24584 9064
rect 24636 9052 24642 9104
rect 24762 9052 24768 9104
rect 24820 9052 24826 9104
rect 25869 9095 25927 9101
rect 25869 9061 25881 9095
rect 25915 9061 25927 9095
rect 25869 9055 25927 9061
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 23952 8928 24225 8956
rect 24213 8925 24225 8928
rect 24259 8925 24271 8959
rect 24213 8919 24271 8925
rect 23569 8891 23627 8897
rect 23569 8857 23581 8891
rect 23615 8888 23627 8891
rect 24780 8888 24808 9052
rect 25884 9024 25912 9055
rect 25700 8996 25912 9024
rect 25521 8959 25579 8965
rect 25521 8925 25533 8959
rect 25567 8956 25579 8959
rect 25700 8956 25728 8996
rect 25567 8928 25728 8956
rect 25777 8959 25835 8965
rect 25567 8925 25579 8928
rect 25521 8919 25579 8925
rect 25777 8925 25789 8959
rect 25823 8925 25835 8959
rect 25976 8956 26004 9132
rect 26050 9120 26056 9172
rect 26108 9120 26114 9172
rect 26068 9024 26096 9120
rect 26068 8996 26372 9024
rect 26344 8965 26372 8996
rect 26053 8959 26111 8965
rect 26053 8956 26065 8959
rect 25976 8928 26065 8956
rect 25777 8919 25835 8925
rect 26053 8925 26065 8928
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26329 8959 26387 8965
rect 26329 8925 26341 8959
rect 26375 8925 26387 8959
rect 26329 8919 26387 8925
rect 23615 8860 24808 8888
rect 23615 8857 23627 8860
rect 23569 8851 23627 8857
rect 25792 8832 25820 8919
rect 22066 8792 22100 8832
rect 22094 8780 22100 8792
rect 22152 8780 22158 8832
rect 23474 8780 23480 8832
rect 23532 8780 23538 8832
rect 24026 8780 24032 8832
rect 24084 8780 24090 8832
rect 25774 8780 25780 8832
rect 25832 8780 25838 8832
rect 25866 8780 25872 8832
rect 25924 8820 25930 8832
rect 26145 8823 26203 8829
rect 26145 8820 26157 8823
rect 25924 8792 26157 8820
rect 25924 8780 25930 8792
rect 26145 8789 26157 8792
rect 26191 8789 26203 8823
rect 26145 8783 26203 8789
rect 1104 8730 31280 8752
rect 1104 8678 4922 8730
rect 4974 8678 4986 8730
rect 5038 8678 5050 8730
rect 5102 8678 5114 8730
rect 5166 8678 5178 8730
rect 5230 8678 5242 8730
rect 5294 8678 10922 8730
rect 10974 8678 10986 8730
rect 11038 8678 11050 8730
rect 11102 8678 11114 8730
rect 11166 8678 11178 8730
rect 11230 8678 11242 8730
rect 11294 8678 16922 8730
rect 16974 8678 16986 8730
rect 17038 8678 17050 8730
rect 17102 8678 17114 8730
rect 17166 8678 17178 8730
rect 17230 8678 17242 8730
rect 17294 8678 22922 8730
rect 22974 8678 22986 8730
rect 23038 8678 23050 8730
rect 23102 8678 23114 8730
rect 23166 8678 23178 8730
rect 23230 8678 23242 8730
rect 23294 8678 28922 8730
rect 28974 8678 28986 8730
rect 29038 8678 29050 8730
rect 29102 8678 29114 8730
rect 29166 8678 29178 8730
rect 29230 8678 29242 8730
rect 29294 8678 31280 8730
rect 1104 8656 31280 8678
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8585 3847 8619
rect 3789 8579 3847 8585
rect 2774 8548 2780 8560
rect 2424 8520 2780 8548
rect 2424 8489 2452 8520
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 3804 8548 3832 8579
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4120 8588 4261 8616
rect 4120 8576 4126 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8576 6058 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7616 8588 7757 8616
rect 7616 8576 7622 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 4614 8548 4620 8560
rect 3804 8520 4620 8548
rect 4614 8508 4620 8520
rect 4672 8548 4678 8560
rect 4985 8551 5043 8557
rect 4985 8548 4997 8551
rect 4672 8520 4997 8548
rect 4672 8508 4678 8520
rect 4985 8517 4997 8520
rect 5031 8517 5043 8551
rect 4985 8511 5043 8517
rect 2682 8489 2688 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2676 8443 2688 8489
rect 2682 8440 2688 8443
rect 2740 8440 2746 8492
rect 3988 8452 4476 8480
rect 3988 8424 4016 8452
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4448 8421 4476 8452
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4856 8452 4905 8480
rect 4856 8440 4862 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5350 8480 5356 8492
rect 5123 8452 5356 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 4341 8415 4399 8421
rect 4341 8412 4353 8415
rect 4120 8384 4353 8412
rect 4120 8372 4126 8384
rect 4341 8381 4353 8384
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 5644 8412 5672 8576
rect 6012 8480 6040 8576
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6012 8452 6377 8480
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6621 8483 6679 8489
rect 6621 8480 6633 8483
rect 6365 8443 6423 8449
rect 6472 8452 6633 8480
rect 6472 8412 6500 8452
rect 6621 8449 6633 8452
rect 6667 8449 6679 8483
rect 7760 8480 7788 8579
rect 7834 8576 7840 8628
rect 7892 8576 7898 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 7984 8588 8984 8616
rect 7984 8576 7990 8588
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 7760 8452 8401 8480
rect 6621 8443 6679 8449
rect 8389 8449 8401 8452
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8662 8480 8668 8492
rect 8619 8452 8668 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8846 8489 8852 8492
rect 8840 8480 8852 8489
rect 8807 8452 8852 8480
rect 8840 8443 8852 8452
rect 8846 8440 8852 8443
rect 8904 8440 8910 8492
rect 8956 8480 8984 8588
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9272 8588 10057 8616
rect 9272 8576 9278 8588
rect 10045 8585 10057 8588
rect 10091 8585 10103 8619
rect 10045 8579 10103 8585
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 11514 8616 11520 8628
rect 10551 8588 11520 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 10413 8483 10471 8489
rect 10413 8480 10425 8483
rect 8956 8452 10425 8480
rect 10413 8449 10425 8452
rect 10459 8480 10471 8483
rect 10502 8480 10508 8492
rect 10459 8452 10508 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 10502 8440 10508 8452
rect 10560 8440 10566 8492
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 11808 8480 11836 8576
rect 11900 8548 11928 8579
rect 12158 8576 12164 8628
rect 12216 8616 12222 8628
rect 12216 8588 12388 8616
rect 12216 8576 12222 8588
rect 12244 8551 12302 8557
rect 12244 8548 12256 8551
rect 11900 8520 12256 8548
rect 12244 8517 12256 8520
rect 12290 8517 12302 8551
rect 12244 8511 12302 8517
rect 11747 8452 11836 8480
rect 11977 8483 12035 8489
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 11977 8449 11989 8483
rect 12023 8480 12035 8483
rect 12360 8480 12388 8588
rect 13354 8576 13360 8628
rect 13412 8576 13418 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8585 15347 8619
rect 15289 8579 15347 8585
rect 12544 8520 14872 8548
rect 12544 8492 12572 8520
rect 12023 8452 12388 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 5644 8384 6500 8412
rect 4433 8375 4491 8381
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 4080 8344 4108 8372
rect 3844 8316 4108 8344
rect 5261 8347 5319 8353
rect 3844 8304 3850 8316
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5307 8316 6408 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 3878 8236 3884 8288
rect 3936 8236 3942 8288
rect 6380 8276 6408 8316
rect 9950 8304 9956 8356
rect 10008 8304 10014 8356
rect 11164 8344 11192 8443
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14844 8489 14872 8520
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 13955 8452 14289 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8480 15255 8483
rect 15304 8480 15332 8579
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15528 8588 15669 8616
rect 15528 8576 15534 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 16485 8619 16543 8625
rect 16485 8585 16497 8619
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 19058 8616 19064 8628
rect 18095 8588 19064 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 16500 8548 16528 8579
rect 16914 8551 16972 8557
rect 16914 8548 16926 8551
rect 16500 8520 16926 8548
rect 16914 8517 16926 8520
rect 16960 8517 16972 8551
rect 16914 8511 16972 8517
rect 15243 8452 15332 8480
rect 15749 8483 15807 8489
rect 15243 8449 15255 8452
rect 15197 8443 15255 8449
rect 15749 8449 15761 8483
rect 15795 8480 15807 8483
rect 16301 8483 16359 8489
rect 15795 8452 16252 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13596 8384 14105 8412
rect 13596 8372 13602 8384
rect 14093 8381 14105 8384
rect 14139 8412 14151 8415
rect 14366 8412 14372 8424
rect 14139 8384 14372 8412
rect 14139 8381 14151 8384
rect 14093 8375 14151 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 16224 8412 16252 8452
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 16574 8480 16580 8492
rect 16347 8452 16580 8480
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 17954 8480 17960 8492
rect 16715 8452 17960 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18524 8489 18552 8588
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19610 8576 19616 8628
rect 19668 8576 19674 8628
rect 19886 8576 19892 8628
rect 19944 8576 19950 8628
rect 20162 8576 20168 8628
rect 20220 8616 20226 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20220 8588 20913 8616
rect 20220 8576 20226 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 21082 8576 21088 8628
rect 21140 8576 21146 8628
rect 21637 8619 21695 8625
rect 21637 8585 21649 8619
rect 21683 8616 21695 8619
rect 21818 8616 21824 8628
rect 21683 8588 21824 8616
rect 21683 8585 21695 8588
rect 21637 8579 21695 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22002 8576 22008 8628
rect 22060 8576 22066 8628
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 23569 8619 23627 8625
rect 23569 8616 23581 8619
rect 23532 8588 23581 8616
rect 23532 8576 23538 8588
rect 23569 8585 23581 8588
rect 23615 8585 23627 8619
rect 23569 8579 23627 8585
rect 24581 8619 24639 8625
rect 24581 8585 24593 8619
rect 24627 8616 24639 8619
rect 24946 8616 24952 8628
rect 24627 8588 24952 8616
rect 24627 8585 24639 8588
rect 24581 8579 24639 8585
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25774 8576 25780 8628
rect 25832 8576 25838 8628
rect 18690 8508 18696 8560
rect 18748 8508 18754 8560
rect 18782 8508 18788 8560
rect 18840 8508 18846 8560
rect 19904 8548 19932 8576
rect 21100 8548 21128 8576
rect 19076 8520 19932 8548
rect 20824 8520 21128 8548
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18598 8440 18604 8492
rect 18656 8440 18662 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8449 18935 8483
rect 18877 8443 18935 8449
rect 16482 8412 16488 8424
rect 16224 8384 16488 8412
rect 15933 8375 15991 8381
rect 13449 8347 13507 8353
rect 13449 8344 13461 8347
rect 11164 8316 12020 8344
rect 7006 8276 7012 8288
rect 6380 8248 7012 8276
rect 7006 8236 7012 8248
rect 7064 8236 7070 8288
rect 11330 8236 11336 8288
rect 11388 8236 11394 8288
rect 11992 8276 12020 8316
rect 12912 8316 13461 8344
rect 12912 8276 12940 8316
rect 13449 8313 13461 8316
rect 13495 8313 13507 8347
rect 15948 8344 15976 8375
rect 16482 8372 16488 8384
rect 16540 8372 16546 8424
rect 18616 8412 18644 8440
rect 18892 8412 18920 8443
rect 18616 8384 18920 8412
rect 16666 8344 16672 8356
rect 15948 8316 16672 8344
rect 13449 8307 13507 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 19076 8353 19104 8520
rect 20824 8489 20852 8520
rect 19705 8483 19763 8489
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 19751 8452 20177 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21453 8483 21511 8489
rect 21453 8449 21465 8483
rect 21499 8480 21511 8483
rect 22020 8480 22048 8576
rect 25792 8548 25820 8576
rect 21499 8452 22048 8480
rect 22112 8520 26004 8548
rect 21499 8449 21511 8452
rect 21453 8443 21511 8449
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8313 19119 8347
rect 19536 8344 19564 8375
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 19812 8344 19840 8372
rect 19536 8316 19840 8344
rect 20073 8347 20131 8353
rect 19061 8307 19119 8313
rect 20073 8313 20085 8347
rect 20119 8344 20131 8347
rect 21100 8344 21128 8443
rect 22112 8424 22140 8520
rect 22364 8483 22422 8489
rect 22364 8449 22376 8483
rect 22410 8480 22422 8483
rect 24026 8480 24032 8492
rect 22410 8452 24032 8480
rect 22410 8449 22422 8452
rect 22364 8443 22422 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 25705 8483 25763 8489
rect 25705 8449 25717 8483
rect 25751 8480 25763 8483
rect 25866 8480 25872 8492
rect 25751 8452 25872 8480
rect 25751 8449 25763 8452
rect 25705 8443 25763 8449
rect 25866 8440 25872 8452
rect 25924 8440 25930 8492
rect 25976 8489 26004 8520
rect 25961 8483 26019 8489
rect 25961 8449 25973 8483
rect 26007 8449 26019 8483
rect 25961 8443 26019 8449
rect 22094 8372 22100 8424
rect 22152 8372 22158 8424
rect 23566 8372 23572 8424
rect 23624 8412 23630 8424
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23624 8384 24133 8412
rect 23624 8372 23630 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 20119 8316 21128 8344
rect 23477 8347 23535 8353
rect 20119 8313 20131 8316
rect 20073 8307 20131 8313
rect 23477 8313 23489 8347
rect 23523 8344 23535 8347
rect 23584 8344 23612 8372
rect 23523 8316 23612 8344
rect 23523 8313 23535 8316
rect 23477 8307 23535 8313
rect 11992 8248 12940 8276
rect 15010 8236 15016 8288
rect 15068 8236 15074 8288
rect 1104 8186 31280 8208
rect 1104 8134 4182 8186
rect 4234 8134 4246 8186
rect 4298 8134 4310 8186
rect 4362 8134 4374 8186
rect 4426 8134 4438 8186
rect 4490 8134 4502 8186
rect 4554 8134 10182 8186
rect 10234 8134 10246 8186
rect 10298 8134 10310 8186
rect 10362 8134 10374 8186
rect 10426 8134 10438 8186
rect 10490 8134 10502 8186
rect 10554 8134 16182 8186
rect 16234 8134 16246 8186
rect 16298 8134 16310 8186
rect 16362 8134 16374 8186
rect 16426 8134 16438 8186
rect 16490 8134 16502 8186
rect 16554 8134 22182 8186
rect 22234 8134 22246 8186
rect 22298 8134 22310 8186
rect 22362 8134 22374 8186
rect 22426 8134 22438 8186
rect 22490 8134 22502 8186
rect 22554 8134 28182 8186
rect 28234 8134 28246 8186
rect 28298 8134 28310 8186
rect 28362 8134 28374 8186
rect 28426 8134 28438 8186
rect 28490 8134 28502 8186
rect 28554 8134 31280 8186
rect 1104 8112 31280 8134
rect 2682 8032 2688 8084
rect 2740 8032 2746 8084
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 7156 8044 7205 8072
rect 7156 8032 7162 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 7193 8035 7251 8041
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12584 8044 12909 8072
rect 12584 8032 12590 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 30742 8032 30748 8084
rect 30800 8032 30806 8084
rect 15930 7964 15936 8016
rect 15988 8004 15994 8016
rect 16117 8007 16175 8013
rect 16117 8004 16129 8007
rect 15988 7976 16129 8004
rect 15988 7964 15994 7976
rect 16117 7973 16129 7976
rect 16163 8004 16175 8007
rect 16163 7976 17816 8004
rect 16163 7973 16175 7976
rect 16117 7967 16175 7973
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7936 16911 7939
rect 17310 7936 17316 7948
rect 16899 7908 17316 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3878 7868 3884 7880
rect 2915 7840 3884 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 9858 7868 9864 7880
rect 6972 7840 9864 7868
rect 6972 7828 6978 7840
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 12158 7868 12164 7880
rect 11563 7840 12164 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7868 14795 7871
rect 14826 7868 14832 7880
rect 14783 7840 14832 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 11348 7800 11376 7828
rect 11762 7803 11820 7809
rect 11762 7800 11774 7803
rect 11348 7772 11774 7800
rect 11762 7769 11774 7772
rect 11808 7769 11820 7803
rect 14476 7800 14504 7831
rect 14826 7828 14832 7840
rect 14884 7828 14890 7880
rect 15010 7877 15016 7880
rect 15004 7868 15016 7877
rect 14971 7840 15016 7868
rect 15004 7831 15016 7840
rect 15010 7828 15016 7831
rect 15068 7828 15074 7880
rect 17788 7877 17816 7976
rect 18322 7964 18328 8016
rect 18380 7964 18386 8016
rect 17589 7871 17647 7877
rect 17589 7868 17601 7871
rect 16316 7840 17601 7868
rect 14476 7772 16252 7800
rect 11762 7763 11820 7769
rect 14642 7692 14648 7744
rect 14700 7692 14706 7744
rect 16224 7741 16252 7772
rect 16316 7744 16344 7840
rect 17589 7837 17601 7840
rect 17635 7837 17647 7871
rect 17589 7831 17647 7837
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17773 7831 17831 7837
rect 17880 7840 18061 7868
rect 16577 7803 16635 7809
rect 16577 7769 16589 7803
rect 16623 7800 16635 7803
rect 17037 7803 17095 7809
rect 17037 7800 17049 7803
rect 16623 7772 17049 7800
rect 16623 7769 16635 7772
rect 16577 7763 16635 7769
rect 17037 7769 17049 7772
rect 17083 7769 17095 7803
rect 17604 7800 17632 7831
rect 17880 7800 17908 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18598 7868 18604 7880
rect 18187 7840 18604 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 30929 7871 30987 7877
rect 30929 7837 30941 7871
rect 30975 7868 30987 7871
rect 31294 7868 31300 7880
rect 30975 7840 31300 7868
rect 30975 7837 30987 7840
rect 30929 7831 30987 7837
rect 31294 7828 31300 7840
rect 31352 7828 31358 7880
rect 17604 7772 17908 7800
rect 17957 7803 18015 7809
rect 17037 7763 17095 7769
rect 17957 7769 17969 7803
rect 18003 7800 18015 7803
rect 18708 7800 18736 7828
rect 18003 7772 18736 7800
rect 18003 7769 18015 7772
rect 17957 7763 18015 7769
rect 16209 7735 16267 7741
rect 16209 7701 16221 7735
rect 16255 7701 16267 7735
rect 16209 7695 16267 7701
rect 16298 7692 16304 7744
rect 16356 7692 16362 7744
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 17862 7732 17868 7744
rect 16724 7704 17868 7732
rect 16724 7692 16730 7704
rect 17862 7692 17868 7704
rect 17920 7732 17926 7744
rect 21634 7732 21640 7744
rect 17920 7704 21640 7732
rect 17920 7692 17926 7704
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 1104 7642 31280 7664
rect 1104 7590 4922 7642
rect 4974 7590 4986 7642
rect 5038 7590 5050 7642
rect 5102 7590 5114 7642
rect 5166 7590 5178 7642
rect 5230 7590 5242 7642
rect 5294 7590 10922 7642
rect 10974 7590 10986 7642
rect 11038 7590 11050 7642
rect 11102 7590 11114 7642
rect 11166 7590 11178 7642
rect 11230 7590 11242 7642
rect 11294 7590 16922 7642
rect 16974 7590 16986 7642
rect 17038 7590 17050 7642
rect 17102 7590 17114 7642
rect 17166 7590 17178 7642
rect 17230 7590 17242 7642
rect 17294 7590 22922 7642
rect 22974 7590 22986 7642
rect 23038 7590 23050 7642
rect 23102 7590 23114 7642
rect 23166 7590 23178 7642
rect 23230 7590 23242 7642
rect 23294 7590 28922 7642
rect 28974 7590 28986 7642
rect 29038 7590 29050 7642
rect 29102 7590 29114 7642
rect 29166 7590 29178 7642
rect 29230 7590 29242 7642
rect 29294 7590 31280 7642
rect 1104 7568 31280 7590
rect 14642 7488 14648 7540
rect 14700 7488 14706 7540
rect 16298 7488 16304 7540
rect 16356 7488 16362 7540
rect 14660 7460 14688 7488
rect 15166 7463 15224 7469
rect 15166 7460 15178 7463
rect 14660 7432 15178 7460
rect 15166 7429 15178 7432
rect 15212 7429 15224 7463
rect 15166 7423 15224 7429
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 14921 7395 14979 7401
rect 14921 7392 14933 7395
rect 14884 7364 14933 7392
rect 14884 7352 14890 7364
rect 14921 7361 14933 7364
rect 14967 7361 14979 7395
rect 14921 7355 14979 7361
rect 1104 7098 31280 7120
rect 1104 7046 4182 7098
rect 4234 7046 4246 7098
rect 4298 7046 4310 7098
rect 4362 7046 4374 7098
rect 4426 7046 4438 7098
rect 4490 7046 4502 7098
rect 4554 7046 10182 7098
rect 10234 7046 10246 7098
rect 10298 7046 10310 7098
rect 10362 7046 10374 7098
rect 10426 7046 10438 7098
rect 10490 7046 10502 7098
rect 10554 7046 16182 7098
rect 16234 7046 16246 7098
rect 16298 7046 16310 7098
rect 16362 7046 16374 7098
rect 16426 7046 16438 7098
rect 16490 7046 16502 7098
rect 16554 7046 22182 7098
rect 22234 7046 22246 7098
rect 22298 7046 22310 7098
rect 22362 7046 22374 7098
rect 22426 7046 22438 7098
rect 22490 7046 22502 7098
rect 22554 7046 28182 7098
rect 28234 7046 28246 7098
rect 28298 7046 28310 7098
rect 28362 7046 28374 7098
rect 28426 7046 28438 7098
rect 28490 7046 28502 7098
rect 28554 7046 31280 7098
rect 1104 7024 31280 7046
rect 20990 6984 20996 6996
rect 18984 6956 20996 6984
rect 5920 6820 6684 6848
rect 5920 6792 5948 6820
rect 5902 6740 5908 6792
rect 5960 6740 5966 6792
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6135 6752 6408 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 6380 6653 6408 6752
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6613 6423 6647
rect 6656 6644 6684 6820
rect 6822 6808 6828 6860
rect 6880 6848 6886 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6880 6820 6929 6848
rect 6880 6808 6886 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 18984 6848 19012 6956
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 22646 6984 22652 6996
rect 21836 6956 22652 6984
rect 19061 6919 19119 6925
rect 19061 6885 19073 6919
rect 19107 6885 19119 6919
rect 19061 6879 19119 6885
rect 19306 6888 21772 6916
rect 7984 6820 8432 6848
rect 7984 6808 7990 6820
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7064 6752 8033 6780
rect 7064 6740 7070 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8404 6789 8432 6820
rect 18708 6820 19012 6848
rect 19076 6848 19104 6879
rect 19306 6848 19334 6888
rect 19076 6820 19334 6848
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8478 6740 8484 6792
rect 8536 6789 8542 6792
rect 8536 6780 8544 6789
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 8536 6752 8581 6780
rect 9692 6752 10517 6780
rect 8536 6743 8544 6752
rect 8536 6740 8542 6743
rect 6733 6715 6791 6721
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 6779 6684 7297 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7285 6681 7297 6684
rect 7331 6681 7343 6715
rect 7285 6675 7343 6681
rect 9692 6656 9720 6752
rect 10505 6749 10517 6752
rect 10551 6780 10563 6783
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10551 6752 10701 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 10689 6749 10701 6752
rect 10735 6749 10747 6783
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10689 6743 10747 6749
rect 10796 6752 10977 6780
rect 10796 6724 10824 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 11422 6780 11428 6792
rect 11103 6752 11428 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 18322 6740 18328 6792
rect 18380 6780 18386 6792
rect 18708 6789 18736 6820
rect 19794 6808 19800 6860
rect 19852 6808 19858 6860
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18380 6752 18429 6780
rect 18380 6740 18386 6752
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 18565 6783 18623 6789
rect 18565 6749 18577 6783
rect 18611 6780 18623 6783
rect 18693 6783 18751 6789
rect 18611 6749 18644 6780
rect 18565 6743 18644 6749
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18923 6783 18981 6789
rect 18923 6749 18935 6783
rect 18969 6780 18981 6783
rect 19426 6780 19432 6792
rect 18969 6752 19432 6780
rect 18969 6749 18981 6752
rect 18923 6743 18981 6749
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6712 10931 6715
rect 11532 6712 11560 6740
rect 10919 6684 11560 6712
rect 10919 6681 10931 6684
rect 10873 6675 10931 6681
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6656 6616 6837 6644
rect 6365 6607 6423 6613
rect 6825 6613 6837 6616
rect 6871 6644 6883 6647
rect 8018 6644 8024 6656
rect 6871 6616 8024 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 9950 6604 9956 6656
rect 10008 6604 10014 6656
rect 11241 6647 11299 6653
rect 11241 6613 11253 6647
rect 11287 6644 11299 6647
rect 11330 6644 11336 6656
rect 11287 6616 11336 6644
rect 11287 6613 11299 6616
rect 11241 6607 11299 6613
rect 11330 6604 11336 6616
rect 11388 6604 11394 6656
rect 18616 6644 18644 6743
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 20714 6780 20720 6792
rect 19536 6752 20720 6780
rect 18785 6715 18843 6721
rect 18785 6681 18797 6715
rect 18831 6712 18843 6715
rect 18831 6684 19380 6712
rect 18831 6681 18843 6684
rect 18785 6675 18843 6681
rect 19150 6644 19156 6656
rect 18616 6616 19156 6644
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19242 6604 19248 6656
rect 19300 6604 19306 6656
rect 19352 6644 19380 6684
rect 19536 6644 19564 6752
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 21085 6783 21143 6789
rect 21085 6749 21097 6783
rect 21131 6780 21143 6783
rect 21131 6752 21220 6780
rect 21131 6749 21143 6752
rect 21085 6743 21143 6749
rect 19613 6715 19671 6721
rect 19613 6681 19625 6715
rect 19659 6712 19671 6715
rect 20073 6715 20131 6721
rect 20073 6712 20085 6715
rect 19659 6684 20085 6712
rect 19659 6681 19671 6684
rect 19613 6675 19671 6681
rect 20073 6681 20085 6684
rect 20119 6681 20131 6715
rect 20073 6675 20131 6681
rect 19352 6616 19564 6644
rect 19702 6604 19708 6656
rect 19760 6604 19766 6656
rect 19794 6604 19800 6656
rect 19852 6644 19858 6656
rect 20806 6644 20812 6656
rect 19852 6616 20812 6644
rect 19852 6604 19858 6616
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 20901 6647 20959 6653
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 20990 6644 20996 6656
rect 20947 6616 20996 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 21192 6653 21220 6752
rect 21634 6740 21640 6792
rect 21692 6740 21698 6792
rect 21744 6780 21772 6888
rect 21836 6857 21864 6956
rect 22646 6944 22652 6956
rect 22704 6944 22710 6996
rect 25133 6987 25191 6993
rect 25133 6953 25145 6987
rect 25179 6953 25191 6987
rect 25133 6947 25191 6953
rect 21821 6851 21879 6857
rect 21821 6817 21833 6851
rect 21867 6817 21879 6851
rect 25148 6848 25176 6947
rect 21821 6811 21879 6817
rect 22112 6820 25176 6848
rect 22112 6780 22140 6820
rect 21744 6752 22140 6780
rect 22189 6783 22247 6789
rect 22189 6749 22201 6783
rect 22235 6749 22247 6783
rect 22189 6743 22247 6749
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 22646 6780 22652 6792
rect 22603 6752 22652 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 22204 6712 22232 6743
rect 22646 6740 22652 6752
rect 22704 6740 22710 6792
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 22756 6752 24409 6780
rect 22020 6684 22232 6712
rect 22373 6715 22431 6721
rect 22020 6656 22048 6684
rect 22373 6681 22385 6715
rect 22419 6681 22431 6715
rect 22373 6675 22431 6681
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 21542 6604 21548 6656
rect 21600 6604 21606 6656
rect 22002 6604 22008 6656
rect 22060 6604 22066 6656
rect 22388 6644 22416 6675
rect 22462 6672 22468 6724
rect 22520 6672 22526 6724
rect 22646 6644 22652 6656
rect 22388 6616 22652 6644
rect 22646 6604 22652 6616
rect 22704 6604 22710 6656
rect 22756 6653 22784 6752
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 24490 6783 24548 6789
rect 24490 6749 24502 6783
rect 24536 6749 24548 6783
rect 24490 6743 24548 6749
rect 24302 6672 24308 6724
rect 24360 6712 24366 6724
rect 24504 6712 24532 6743
rect 24578 6740 24584 6792
rect 24636 6780 24642 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24636 6752 24685 6780
rect 24636 6740 24642 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 24854 6740 24860 6792
rect 24912 6789 24918 6792
rect 24912 6743 24920 6789
rect 24912 6740 24918 6743
rect 25130 6740 25136 6792
rect 25188 6740 25194 6792
rect 25225 6783 25283 6789
rect 25225 6749 25237 6783
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 24360 6684 24532 6712
rect 24360 6672 24366 6684
rect 24762 6672 24768 6724
rect 24820 6672 24826 6724
rect 25240 6712 25268 6743
rect 25056 6684 25268 6712
rect 25056 6653 25084 6684
rect 22741 6647 22799 6653
rect 22741 6613 22753 6647
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 25041 6647 25099 6653
rect 25041 6613 25053 6647
rect 25087 6613 25099 6647
rect 25041 6607 25099 6613
rect 25501 6647 25559 6653
rect 25501 6613 25513 6647
rect 25547 6644 25559 6647
rect 26234 6644 26240 6656
rect 25547 6616 26240 6644
rect 25547 6613 25559 6616
rect 25501 6607 25559 6613
rect 26234 6604 26240 6616
rect 26292 6604 26298 6656
rect 1104 6554 31280 6576
rect 1104 6502 4922 6554
rect 4974 6502 4986 6554
rect 5038 6502 5050 6554
rect 5102 6502 5114 6554
rect 5166 6502 5178 6554
rect 5230 6502 5242 6554
rect 5294 6502 10922 6554
rect 10974 6502 10986 6554
rect 11038 6502 11050 6554
rect 11102 6502 11114 6554
rect 11166 6502 11178 6554
rect 11230 6502 11242 6554
rect 11294 6502 16922 6554
rect 16974 6502 16986 6554
rect 17038 6502 17050 6554
rect 17102 6502 17114 6554
rect 17166 6502 17178 6554
rect 17230 6502 17242 6554
rect 17294 6502 22922 6554
rect 22974 6502 22986 6554
rect 23038 6502 23050 6554
rect 23102 6502 23114 6554
rect 23166 6502 23178 6554
rect 23230 6502 23242 6554
rect 23294 6502 28922 6554
rect 28974 6502 28986 6554
rect 29038 6502 29050 6554
rect 29102 6502 29114 6554
rect 29166 6502 29178 6554
rect 29230 6502 29242 6554
rect 29294 6502 31280 6554
rect 1104 6480 31280 6502
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5460 6304 5488 6403
rect 5902 6400 5908 6452
rect 5960 6400 5966 6452
rect 5994 6400 6000 6452
rect 6052 6400 6058 6452
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6440 7803 6443
rect 7926 6440 7932 6452
rect 7791 6412 7932 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8018 6400 8024 6452
rect 8076 6400 8082 6452
rect 8662 6400 8668 6452
rect 8720 6400 8726 6452
rect 9674 6400 9680 6452
rect 9732 6400 9738 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 10008 6412 10149 6440
rect 10008 6400 10014 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14093 6443 14151 6449
rect 14093 6440 14105 6443
rect 13872 6412 14105 6440
rect 13872 6400 13878 6412
rect 14093 6409 14105 6412
rect 14139 6409 14151 6443
rect 14093 6403 14151 6409
rect 19242 6400 19248 6452
rect 19300 6400 19306 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 20772 6412 20821 6440
rect 20772 6400 20778 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 21542 6400 21548 6452
rect 21600 6440 21606 6452
rect 21913 6443 21971 6449
rect 21913 6440 21925 6443
rect 21600 6412 21925 6440
rect 21600 6400 21606 6412
rect 21913 6409 21925 6412
rect 21959 6409 21971 6443
rect 21913 6403 21971 6409
rect 22462 6400 22468 6452
rect 22520 6400 22526 6452
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 23753 6443 23811 6449
rect 23753 6440 23765 6443
rect 23624 6412 23765 6440
rect 23624 6400 23630 6412
rect 23753 6409 23765 6412
rect 23799 6440 23811 6443
rect 24210 6440 24216 6452
rect 23799 6412 24216 6440
rect 23799 6409 23811 6412
rect 23753 6403 23811 6409
rect 24210 6400 24216 6412
rect 24268 6440 24274 6452
rect 24581 6443 24639 6449
rect 24581 6440 24593 6443
rect 24268 6412 24593 6440
rect 24268 6400 24274 6412
rect 24581 6409 24593 6412
rect 24627 6440 24639 6443
rect 24670 6440 24676 6452
rect 24627 6412 24676 6440
rect 24627 6409 24639 6412
rect 24581 6403 24639 6409
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 24762 6400 24768 6452
rect 24820 6440 24826 6452
rect 24820 6412 26372 6440
rect 24820 6400 24826 6412
rect 5215 6276 5488 6304
rect 5813 6307 5871 6313
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 6012 6304 6040 6400
rect 8680 6372 8708 6400
rect 19260 6372 19288 6400
rect 22094 6372 22100 6384
rect 6380 6344 8340 6372
rect 8680 6344 10732 6372
rect 6380 6313 6408 6344
rect 8312 6313 8340 6344
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6012 6276 6377 6304
rect 5813 6267 5871 6273
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6621 6307 6679 6313
rect 6621 6304 6633 6307
rect 6365 6267 6423 6273
rect 6472 6276 6633 6304
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 5828 6168 5856 6267
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6178 6236 6184 6248
rect 6135 6208 6184 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6472 6236 6500 6276
rect 6621 6273 6633 6276
rect 6667 6273 6679 6307
rect 6621 6267 6679 6273
rect 7837 6307 7895 6313
rect 7837 6273 7849 6307
rect 7883 6304 7895 6307
rect 8297 6307 8355 6313
rect 7883 6276 8156 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 6328 6208 6500 6236
rect 6328 6196 6334 6208
rect 6362 6168 6368 6180
rect 4120 6140 5488 6168
rect 5828 6140 6368 6168
rect 4120 6128 4126 6140
rect 5350 6060 5356 6112
rect 5408 6060 5414 6112
rect 5460 6100 5488 6140
rect 6362 6128 6368 6140
rect 6420 6128 6426 6180
rect 8128 6168 8156 6276
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8564 6307 8622 6313
rect 8564 6273 8576 6307
rect 8610 6304 8622 6307
rect 8938 6304 8944 6316
rect 8610 6276 8944 6304
rect 8610 6273 8622 6276
rect 8564 6267 8622 6273
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10100 6276 10364 6304
rect 10100 6264 10106 6276
rect 10336 6245 10364 6276
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6205 10379 6239
rect 10321 6199 10379 6205
rect 10244 6168 10272 6199
rect 7300 6140 8156 6168
rect 7300 6100 7328 6140
rect 5460 6072 7328 6100
rect 8128 6100 8156 6140
rect 9232 6140 10272 6168
rect 9232 6100 9260 6140
rect 8128 6072 9260 6100
rect 9766 6060 9772 6112
rect 9824 6060 9830 6112
rect 10594 6060 10600 6112
rect 10652 6060 10658 6112
rect 10704 6100 10732 6344
rect 17696 6344 19288 6372
rect 19444 6344 22100 6372
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11974 6304 11980 6316
rect 11563 6276 11980 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 17696 6313 17724 6344
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 14185 6307 14243 6313
rect 13495 6276 13768 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 10836 6208 11161 6236
rect 10836 6196 10842 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 11606 6196 11612 6248
rect 11664 6196 11670 6248
rect 13740 6177 13768 6276
rect 14185 6273 14197 6307
rect 14231 6304 14243 6307
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 14231 6276 14565 6304
rect 14231 6273 14243 6276
rect 14185 6267 14243 6273
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 17954 6264 17960 6316
rect 18012 6264 18018 6316
rect 18230 6313 18236 6316
rect 18224 6267 18236 6313
rect 18230 6264 18236 6267
rect 18288 6264 18294 6316
rect 19444 6313 19472 6344
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19685 6307 19743 6313
rect 19685 6304 19697 6307
rect 19429 6267 19487 6273
rect 19536 6276 19697 6304
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 13872 6208 14289 6236
rect 13872 6196 13878 6208
rect 14200 6180 14228 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 15194 6196 15200 6248
rect 15252 6196 15258 6248
rect 19536 6236 19564 6276
rect 19685 6273 19697 6276
rect 19731 6273 19743 6307
rect 22480 6304 22508 6400
rect 23661 6375 23719 6381
rect 23661 6341 23673 6375
rect 23707 6372 23719 6375
rect 25041 6375 25099 6381
rect 25041 6372 25053 6375
rect 23707 6344 25053 6372
rect 23707 6341 23719 6344
rect 23661 6335 23719 6341
rect 25041 6341 25053 6344
rect 25087 6341 25099 6375
rect 25041 6335 25099 6341
rect 23198 6304 23204 6316
rect 22480 6276 23204 6304
rect 19685 6267 19743 6273
rect 23198 6264 23204 6276
rect 23256 6264 23262 6316
rect 24394 6264 24400 6316
rect 24452 6304 24458 6316
rect 26344 6313 26372 6412
rect 24673 6307 24731 6313
rect 24452 6276 24624 6304
rect 24452 6264 24458 6276
rect 19260 6208 19564 6236
rect 21453 6239 21511 6245
rect 13725 6171 13783 6177
rect 13725 6137 13737 6171
rect 13771 6137 13783 6171
rect 13725 6131 13783 6137
rect 14182 6128 14188 6180
rect 14240 6128 14246 6180
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 10704 6072 11529 6100
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 11882 6060 11888 6112
rect 11940 6060 11946 6112
rect 13630 6060 13636 6112
rect 13688 6060 13694 6112
rect 17865 6103 17923 6109
rect 17865 6069 17877 6103
rect 17911 6100 17923 6103
rect 19260 6100 19288 6208
rect 21453 6205 21465 6239
rect 21499 6205 21511 6239
rect 21453 6199 21511 6205
rect 20438 6128 20444 6180
rect 20496 6168 20502 6180
rect 20901 6171 20959 6177
rect 20901 6168 20913 6171
rect 20496 6140 20913 6168
rect 20496 6128 20502 6140
rect 20901 6137 20913 6140
rect 20947 6137 20959 6171
rect 20901 6131 20959 6137
rect 17911 6072 19288 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 19334 6060 19340 6112
rect 19392 6100 19398 6112
rect 21468 6100 21496 6199
rect 22002 6196 22008 6248
rect 22060 6236 22066 6248
rect 22465 6239 22523 6245
rect 22465 6236 22477 6239
rect 22060 6208 22477 6236
rect 22060 6196 22066 6208
rect 22465 6205 22477 6208
rect 22511 6205 22523 6239
rect 22465 6199 22523 6205
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6236 23627 6239
rect 24596 6236 24624 6276
rect 24673 6273 24685 6307
rect 24719 6304 24731 6307
rect 25777 6307 25835 6313
rect 25777 6304 25789 6307
rect 24719 6276 25789 6304
rect 24719 6273 24731 6276
rect 24673 6267 24731 6273
rect 25777 6273 25789 6276
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 26329 6307 26387 6313
rect 26329 6273 26341 6307
rect 26375 6273 26387 6307
rect 26329 6267 26387 6273
rect 24765 6239 24823 6245
rect 24765 6236 24777 6239
rect 23615 6208 24532 6236
rect 24596 6208 24777 6236
rect 23615 6205 23627 6208
rect 23569 6199 23627 6205
rect 24302 6128 24308 6180
rect 24360 6128 24366 6180
rect 24504 6168 24532 6208
rect 24765 6205 24777 6208
rect 24811 6205 24823 6239
rect 25593 6239 25651 6245
rect 25593 6236 25605 6239
rect 24765 6199 24823 6205
rect 25516 6208 25605 6236
rect 25406 6168 25412 6180
rect 24504 6140 25412 6168
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 19392 6072 21496 6100
rect 19392 6060 19398 6072
rect 22646 6060 22652 6112
rect 22704 6060 22710 6112
rect 24118 6060 24124 6112
rect 24176 6060 24182 6112
rect 24210 6060 24216 6112
rect 24268 6060 24274 6112
rect 24320 6100 24348 6128
rect 25516 6100 25544 6208
rect 25593 6205 25605 6208
rect 25639 6205 25651 6239
rect 25593 6199 25651 6205
rect 24320 6072 25544 6100
rect 1104 6010 31280 6032
rect 1104 5958 4182 6010
rect 4234 5958 4246 6010
rect 4298 5958 4310 6010
rect 4362 5958 4374 6010
rect 4426 5958 4438 6010
rect 4490 5958 4502 6010
rect 4554 5958 10182 6010
rect 10234 5958 10246 6010
rect 10298 5958 10310 6010
rect 10362 5958 10374 6010
rect 10426 5958 10438 6010
rect 10490 5958 10502 6010
rect 10554 5958 16182 6010
rect 16234 5958 16246 6010
rect 16298 5958 16310 6010
rect 16362 5958 16374 6010
rect 16426 5958 16438 6010
rect 16490 5958 16502 6010
rect 16554 5958 22182 6010
rect 22234 5958 22246 6010
rect 22298 5958 22310 6010
rect 22362 5958 22374 6010
rect 22426 5958 22438 6010
rect 22490 5958 22502 6010
rect 22554 5958 28182 6010
rect 28234 5958 28246 6010
rect 28298 5958 28310 6010
rect 28362 5958 28374 6010
rect 28426 5958 28438 6010
rect 28490 5958 28502 6010
rect 28554 5958 31280 6010
rect 1104 5936 31280 5958
rect 5350 5856 5356 5908
rect 5408 5856 5414 5908
rect 5994 5896 6000 5908
rect 5644 5868 6000 5896
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 5368 5692 5396 5856
rect 5644 5769 5672 5868
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6420 5868 7113 5896
rect 6420 5856 6426 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 7101 5859 7159 5865
rect 8110 5856 8116 5908
rect 8168 5856 8174 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 9766 5856 9772 5908
rect 9824 5856 9830 5908
rect 10594 5896 10600 5908
rect 10152 5868 10600 5896
rect 7009 5831 7067 5837
rect 7009 5797 7021 5831
rect 7055 5828 7067 5831
rect 7055 5800 7788 5828
rect 7055 5797 7067 5800
rect 7009 5791 7067 5797
rect 7760 5769 7788 5800
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8128 5760 8156 5856
rect 7791 5732 8156 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 5885 5695 5943 5701
rect 5885 5692 5897 5695
rect 5368 5664 5897 5692
rect 5885 5661 5897 5664
rect 5931 5661 5943 5695
rect 5885 5655 5943 5661
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9784 5692 9812 5856
rect 10152 5769 10180 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 11664 5868 11989 5896
rect 11664 5856 11670 5868
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 13630 5856 13636 5908
rect 13688 5856 13694 5908
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15252 5868 15485 5896
rect 15252 5856 15258 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 18230 5856 18236 5908
rect 18288 5896 18294 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 18288 5868 18337 5896
rect 18288 5856 18294 5868
rect 18325 5865 18337 5868
rect 18371 5865 18383 5899
rect 18325 5859 18383 5865
rect 20732 5868 21772 5896
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10686 5760 10692 5772
rect 10367 5732 10692 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 13538 5760 13544 5772
rect 11195 5732 13544 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 9171 5664 9812 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 11330 5652 11336 5704
rect 11388 5652 11394 5704
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 11480 5664 11525 5692
rect 11480 5652 11486 5664
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 11839 5695 11897 5701
rect 11839 5661 11851 5695
rect 11885 5692 11897 5695
rect 12066 5692 12072 5704
rect 11885 5664 12072 5692
rect 11885 5661 11897 5664
rect 11839 5655 11897 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 8036 5624 8064 5652
rect 10045 5627 10103 5633
rect 10045 5624 10057 5627
rect 8036 5596 10057 5624
rect 10045 5593 10057 5596
rect 10091 5624 10103 5627
rect 10594 5624 10600 5636
rect 10091 5596 10600 5624
rect 10091 5593 10103 5596
rect 10045 5587 10103 5593
rect 10594 5584 10600 5596
rect 10652 5624 10658 5636
rect 10873 5627 10931 5633
rect 10873 5624 10885 5627
rect 10652 5596 10885 5624
rect 10652 5584 10658 5596
rect 10873 5593 10885 5596
rect 10919 5593 10931 5627
rect 10873 5587 10931 5593
rect 11698 5584 11704 5636
rect 11756 5584 11762 5636
rect 13648 5624 13676 5856
rect 20438 5788 20444 5840
rect 20496 5788 20502 5840
rect 19889 5763 19947 5769
rect 19889 5729 19901 5763
rect 19935 5760 19947 5763
rect 19978 5760 19984 5772
rect 19935 5732 19984 5760
rect 19935 5729 19947 5732
rect 19889 5723 19947 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14826 5692 14832 5704
rect 14139 5664 14832 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 19613 5695 19671 5701
rect 18555 5664 19288 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 14338 5627 14396 5633
rect 14338 5624 14350 5627
rect 13648 5596 14350 5624
rect 14338 5593 14350 5596
rect 14384 5593 14396 5627
rect 14338 5587 14396 5593
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 4062 5556 4068 5568
rect 1627 5528 4068 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 4062 5516 4068 5528
rect 4120 5516 4126 5568
rect 9674 5516 9680 5568
rect 9732 5516 9738 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 10192 5528 10517 5556
rect 10192 5516 10198 5528
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 10505 5519 10563 5525
rect 10965 5559 11023 5565
rect 10965 5525 10977 5559
rect 11011 5556 11023 5559
rect 11514 5556 11520 5568
rect 11011 5528 11520 5556
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 19260 5565 19288 5664
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 20456 5692 20484 5788
rect 20732 5701 20760 5868
rect 20990 5701 20996 5704
rect 19659 5664 20484 5692
rect 20717 5695 20775 5701
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 20717 5661 20729 5695
rect 20763 5661 20775 5695
rect 20717 5655 20775 5661
rect 20984 5655 20996 5701
rect 21048 5692 21054 5704
rect 21744 5692 21772 5868
rect 22002 5856 22008 5908
rect 22060 5896 22066 5908
rect 22097 5899 22155 5905
rect 22097 5896 22109 5899
rect 22060 5868 22109 5896
rect 22060 5856 22066 5868
rect 22097 5865 22109 5868
rect 22143 5865 22155 5899
rect 22097 5859 22155 5865
rect 23198 5856 23204 5908
rect 23256 5896 23262 5908
rect 23569 5899 23627 5905
rect 23569 5896 23581 5899
rect 23256 5868 23581 5896
rect 23256 5856 23262 5868
rect 23569 5865 23581 5868
rect 23615 5865 23627 5899
rect 23569 5859 23627 5865
rect 24118 5856 24124 5908
rect 24176 5856 24182 5908
rect 24210 5856 24216 5908
rect 24268 5856 24274 5908
rect 24762 5856 24768 5908
rect 24820 5896 24826 5908
rect 25777 5899 25835 5905
rect 25777 5896 25789 5899
rect 24820 5868 25789 5896
rect 24820 5856 24826 5868
rect 25777 5865 25789 5868
rect 25823 5865 25835 5899
rect 25777 5859 25835 5865
rect 24136 5760 24164 5856
rect 23860 5732 24164 5760
rect 22094 5692 22100 5704
rect 21048 5664 21084 5692
rect 21744 5664 22100 5692
rect 20990 5652 20996 5655
rect 21048 5652 21054 5664
rect 22094 5652 22100 5664
rect 22152 5692 22158 5704
rect 23860 5701 23888 5732
rect 22189 5695 22247 5701
rect 22189 5692 22201 5695
rect 22152 5664 22201 5692
rect 22152 5652 22158 5664
rect 22189 5661 22201 5664
rect 22235 5692 22247 5695
rect 23845 5695 23903 5701
rect 22235 5664 23428 5692
rect 22235 5661 22247 5664
rect 22189 5655 22247 5661
rect 23400 5636 23428 5664
rect 23845 5661 23857 5695
rect 23891 5661 23903 5695
rect 23845 5655 23903 5661
rect 23937 5695 23995 5701
rect 23937 5661 23949 5695
rect 23983 5692 23995 5695
rect 24228 5692 24256 5856
rect 25406 5788 25412 5840
rect 25464 5828 25470 5840
rect 25869 5831 25927 5837
rect 25869 5828 25881 5831
rect 25464 5800 25881 5828
rect 25464 5788 25470 5800
rect 25869 5797 25881 5800
rect 25915 5797 25927 5831
rect 25869 5791 25927 5797
rect 26510 5720 26516 5772
rect 26568 5720 26574 5772
rect 23983 5664 24256 5692
rect 24397 5695 24455 5701
rect 23983 5661 23995 5664
rect 23937 5655 23995 5661
rect 24397 5661 24409 5695
rect 24443 5692 24455 5695
rect 25498 5692 25504 5704
rect 24443 5664 25504 5692
rect 24443 5661 24455 5664
rect 24397 5655 24455 5661
rect 22278 5584 22284 5636
rect 22336 5624 22342 5636
rect 22434 5627 22492 5633
rect 22434 5624 22446 5627
rect 22336 5596 22446 5624
rect 22336 5584 22342 5596
rect 22434 5593 22446 5596
rect 22480 5593 22492 5627
rect 22434 5587 22492 5593
rect 23382 5584 23388 5636
rect 23440 5624 23446 5636
rect 24412 5624 24440 5655
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 26237 5695 26295 5701
rect 26237 5661 26249 5695
rect 26283 5661 26295 5695
rect 26237 5655 26295 5661
rect 24642 5627 24700 5633
rect 24642 5624 24654 5627
rect 23440 5596 24440 5624
rect 24504 5596 24654 5624
rect 23440 5584 23446 5596
rect 19245 5559 19303 5565
rect 19245 5525 19257 5559
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 19702 5516 19708 5568
rect 19760 5556 19766 5568
rect 22186 5556 22192 5568
rect 19760 5528 22192 5556
rect 19760 5516 19766 5528
rect 22186 5516 22192 5528
rect 22244 5556 22250 5568
rect 23566 5556 23572 5568
rect 22244 5528 23572 5556
rect 22244 5516 22250 5528
rect 23566 5516 23572 5528
rect 23624 5516 23630 5568
rect 23658 5516 23664 5568
rect 23716 5516 23722 5568
rect 24121 5559 24179 5565
rect 24121 5525 24133 5559
rect 24167 5556 24179 5559
rect 24504 5556 24532 5596
rect 24642 5593 24654 5596
rect 24688 5593 24700 5627
rect 24642 5587 24700 5593
rect 24762 5584 24768 5636
rect 24820 5624 24826 5636
rect 26252 5624 26280 5655
rect 27062 5652 27068 5704
rect 27120 5692 27126 5704
rect 27249 5695 27307 5701
rect 27249 5692 27261 5695
rect 27120 5664 27261 5692
rect 27120 5652 27126 5664
rect 27249 5661 27261 5664
rect 27295 5661 27307 5695
rect 27249 5655 27307 5661
rect 24820 5596 26280 5624
rect 24820 5584 24826 5596
rect 24167 5528 24532 5556
rect 26329 5559 26387 5565
rect 24167 5525 24179 5528
rect 24121 5519 24179 5525
rect 26329 5525 26341 5559
rect 26375 5556 26387 5559
rect 26697 5559 26755 5565
rect 26697 5556 26709 5559
rect 26375 5528 26709 5556
rect 26375 5525 26387 5528
rect 26329 5519 26387 5525
rect 26697 5525 26709 5528
rect 26743 5525 26755 5559
rect 26697 5519 26755 5525
rect 1104 5466 31280 5488
rect 1104 5414 4922 5466
rect 4974 5414 4986 5466
rect 5038 5414 5050 5466
rect 5102 5414 5114 5466
rect 5166 5414 5178 5466
rect 5230 5414 5242 5466
rect 5294 5414 10922 5466
rect 10974 5414 10986 5466
rect 11038 5414 11050 5466
rect 11102 5414 11114 5466
rect 11166 5414 11178 5466
rect 11230 5414 11242 5466
rect 11294 5414 16922 5466
rect 16974 5414 16986 5466
rect 17038 5414 17050 5466
rect 17102 5414 17114 5466
rect 17166 5414 17178 5466
rect 17230 5414 17242 5466
rect 17294 5414 22922 5466
rect 22974 5414 22986 5466
rect 23038 5414 23050 5466
rect 23102 5414 23114 5466
rect 23166 5414 23178 5466
rect 23230 5414 23242 5466
rect 23294 5414 28922 5466
rect 28974 5414 28986 5466
rect 29038 5414 29050 5466
rect 29102 5414 29114 5466
rect 29166 5414 29178 5466
rect 29230 5414 29242 5466
rect 29294 5414 31280 5466
rect 1104 5392 31280 5414
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 10778 5352 10784 5364
rect 10643 5324 10784 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 12676 5324 12940 5352
rect 12676 5312 12682 5324
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12342 5284 12348 5296
rect 12124 5256 12348 5284
rect 12124 5244 12130 5256
rect 12342 5244 12348 5256
rect 12400 5284 12406 5296
rect 12912 5293 12940 5324
rect 15286 5312 15292 5364
rect 15344 5312 15350 5364
rect 21821 5355 21879 5361
rect 21821 5321 21833 5355
rect 21867 5321 21879 5355
rect 21821 5315 21879 5321
rect 12897 5287 12955 5293
rect 12400 5256 12848 5284
rect 12400 5244 12406 5256
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 9214 5216 9220 5228
rect 8812 5188 9220 5216
rect 8812 5176 8818 5188
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9306 5176 9312 5228
rect 9364 5216 9370 5228
rect 9473 5219 9531 5225
rect 9473 5216 9485 5219
rect 9364 5188 9485 5216
rect 9364 5176 9370 5188
rect 9473 5185 9485 5188
rect 9519 5185 9531 5219
rect 9473 5179 9531 5185
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12820 5216 12848 5256
rect 12897 5253 12909 5287
rect 12943 5253 12955 5287
rect 12897 5247 12955 5253
rect 12989 5287 13047 5293
rect 12989 5253 13001 5287
rect 13035 5284 13047 5287
rect 13357 5287 13415 5293
rect 13357 5284 13369 5287
rect 13035 5256 13369 5284
rect 13035 5253 13047 5256
rect 12989 5247 13047 5253
rect 13357 5253 13369 5256
rect 13403 5253 13415 5287
rect 15304 5284 15332 5312
rect 17770 5284 17776 5296
rect 13357 5247 13415 5253
rect 15028 5256 17776 5284
rect 15028 5225 15056 5256
rect 17770 5244 17776 5256
rect 17828 5244 17834 5296
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12820 5188 13093 5216
rect 12713 5179 12771 5185
rect 13081 5185 13093 5188
rect 13127 5216 13139 5219
rect 15013 5219 15071 5225
rect 13127 5188 14780 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 11422 5108 11428 5160
rect 11480 5148 11486 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11480 5120 12081 5148
rect 11480 5108 11486 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 12728 5080 12756 5179
rect 13906 5108 13912 5160
rect 13964 5108 13970 5160
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14645 5151 14703 5157
rect 14645 5148 14657 5151
rect 14424 5120 14657 5148
rect 14424 5108 14430 5120
rect 14645 5117 14657 5120
rect 14691 5117 14703 5151
rect 14752 5148 14780 5188
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 15289 5219 15347 5225
rect 15289 5216 15301 5219
rect 15252 5188 15301 5216
rect 15252 5176 15258 5188
rect 15289 5185 15301 5188
rect 15335 5185 15347 5219
rect 15289 5179 15347 5185
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5216 21235 5219
rect 21836 5216 21864 5315
rect 22186 5312 22192 5364
rect 22244 5312 22250 5364
rect 22281 5355 22339 5361
rect 22281 5321 22293 5355
rect 22327 5352 22339 5355
rect 22646 5352 22652 5364
rect 22327 5324 22652 5352
rect 22327 5321 22339 5324
rect 22281 5315 22339 5321
rect 22646 5312 22652 5324
rect 22704 5312 22710 5364
rect 23382 5312 23388 5364
rect 23440 5312 23446 5364
rect 24302 5312 24308 5364
rect 24360 5312 24366 5364
rect 25317 5355 25375 5361
rect 25317 5321 25329 5355
rect 25363 5321 25375 5355
rect 25317 5315 25375 5321
rect 23400 5284 23428 5312
rect 22940 5256 23428 5284
rect 22940 5225 22968 5256
rect 23658 5244 23664 5296
rect 23716 5244 23722 5296
rect 25332 5284 25360 5315
rect 25654 5287 25712 5293
rect 25654 5284 25666 5287
rect 25332 5256 25666 5284
rect 25654 5253 25666 5256
rect 25700 5253 25712 5287
rect 25654 5247 25712 5253
rect 21223 5188 21864 5216
rect 22925 5219 22983 5225
rect 21223 5185 21235 5188
rect 21177 5179 21235 5185
rect 22925 5185 22937 5219
rect 22971 5185 22983 5219
rect 22925 5179 22983 5185
rect 23192 5219 23250 5225
rect 23192 5185 23204 5219
rect 23238 5216 23250 5219
rect 23676 5216 23704 5244
rect 23238 5188 23704 5216
rect 25133 5219 25191 5225
rect 23238 5185 23250 5188
rect 23192 5179 23250 5185
rect 25133 5185 25145 5219
rect 25179 5216 25191 5219
rect 25314 5216 25320 5228
rect 25179 5188 25320 5216
rect 25179 5185 25191 5188
rect 25133 5179 25191 5185
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 25409 5219 25467 5225
rect 25409 5185 25421 5219
rect 25455 5216 25467 5219
rect 25498 5216 25504 5228
rect 25455 5188 25504 5216
rect 25455 5185 25467 5188
rect 25409 5179 25467 5185
rect 25498 5176 25504 5188
rect 25556 5176 25562 5228
rect 26694 5176 26700 5228
rect 26752 5216 26758 5228
rect 27249 5219 27307 5225
rect 27249 5216 27261 5219
rect 26752 5188 27261 5216
rect 26752 5176 26758 5188
rect 27249 5185 27261 5188
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 22465 5151 22523 5157
rect 14752 5120 17448 5148
rect 14645 5111 14703 5117
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 12728 5052 14841 5080
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 14918 5040 14924 5092
rect 14976 5080 14982 5092
rect 15197 5083 15255 5089
rect 15197 5080 15209 5083
rect 14976 5052 15209 5080
rect 14976 5040 14982 5052
rect 15197 5049 15209 5052
rect 15243 5049 15255 5083
rect 15197 5043 15255 5049
rect 17420 5024 17448 5120
rect 22465 5117 22477 5151
rect 22511 5148 22523 5151
rect 22830 5148 22836 5160
rect 22511 5120 22836 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 22830 5108 22836 5120
rect 22888 5108 22894 5160
rect 26973 5151 27031 5157
rect 26973 5117 26985 5151
rect 27019 5148 27031 5151
rect 27062 5148 27068 5160
rect 27019 5120 27068 5148
rect 27019 5117 27031 5120
rect 26973 5111 27031 5117
rect 21361 5083 21419 5089
rect 21361 5049 21373 5083
rect 21407 5080 21419 5083
rect 22278 5080 22284 5092
rect 21407 5052 22284 5080
rect 21407 5049 21419 5052
rect 21361 5043 21419 5049
rect 22278 5040 22284 5052
rect 22336 5040 22342 5092
rect 26789 5083 26847 5089
rect 26789 5049 26801 5083
rect 26835 5080 26847 5083
rect 26988 5080 27016 5111
rect 27062 5108 27068 5120
rect 27120 5108 27126 5160
rect 26835 5052 27016 5080
rect 26835 5049 26847 5052
rect 26789 5043 26847 5049
rect 12434 4972 12440 5024
rect 12492 4972 12498 5024
rect 13265 5015 13323 5021
rect 13265 4981 13277 5015
rect 13311 5012 13323 5015
rect 13814 5012 13820 5024
rect 13311 4984 13820 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14090 4972 14096 5024
rect 14148 4972 14154 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 16574 5012 16580 5024
rect 14240 4984 16580 5012
rect 14240 4972 14246 4984
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17402 4972 17408 5024
rect 17460 4972 17466 5024
rect 26602 4972 26608 5024
rect 26660 5012 26666 5024
rect 27065 5015 27123 5021
rect 27065 5012 27077 5015
rect 26660 4984 27077 5012
rect 26660 4972 26666 4984
rect 27065 4981 27077 4984
rect 27111 4981 27123 5015
rect 27065 4975 27123 4981
rect 27430 4972 27436 5024
rect 27488 4972 27494 5024
rect 1104 4922 31280 4944
rect 1104 4870 4182 4922
rect 4234 4870 4246 4922
rect 4298 4870 4310 4922
rect 4362 4870 4374 4922
rect 4426 4870 4438 4922
rect 4490 4870 4502 4922
rect 4554 4870 10182 4922
rect 10234 4870 10246 4922
rect 10298 4870 10310 4922
rect 10362 4870 10374 4922
rect 10426 4870 10438 4922
rect 10490 4870 10502 4922
rect 10554 4870 16182 4922
rect 16234 4870 16246 4922
rect 16298 4870 16310 4922
rect 16362 4870 16374 4922
rect 16426 4870 16438 4922
rect 16490 4870 16502 4922
rect 16554 4870 22182 4922
rect 22234 4870 22246 4922
rect 22298 4870 22310 4922
rect 22362 4870 22374 4922
rect 22426 4870 22438 4922
rect 22490 4870 22502 4922
rect 22554 4870 28182 4922
rect 28234 4870 28246 4922
rect 28298 4870 28310 4922
rect 28362 4870 28374 4922
rect 28426 4870 28438 4922
rect 28490 4870 28502 4922
rect 28554 4870 31280 4922
rect 1104 4848 31280 4870
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9364 4780 9505 4808
rect 9364 4768 9370 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 10612 4780 12572 4808
rect 9401 4743 9459 4749
rect 9401 4709 9413 4743
rect 9447 4740 9459 4743
rect 9766 4740 9772 4752
rect 9447 4712 9772 4740
rect 9447 4709 9459 4712
rect 9401 4703 9459 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 10045 4743 10103 4749
rect 10045 4709 10057 4743
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 10060 4672 10088 4703
rect 9232 4644 10088 4672
rect 9232 4613 9260 4644
rect 10612 4616 10640 4780
rect 12253 4743 12311 4749
rect 12253 4709 12265 4743
rect 12299 4709 12311 4743
rect 12544 4740 12572 4780
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12676 4780 13093 4808
rect 12676 4768 12682 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 14090 4808 14096 4820
rect 13081 4771 13139 4777
rect 13556 4780 14096 4808
rect 12544 4712 13492 4740
rect 12253 4703 12311 4709
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 12268 4672 12296 4703
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 10735 4644 11560 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 10042 4604 10048 4616
rect 9999 4576 10048 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 10413 4607 10471 4613
rect 10413 4573 10425 4607
rect 10459 4604 10471 4607
rect 10594 4604 10600 4616
rect 10459 4576 10600 4604
rect 10459 4573 10471 4576
rect 10413 4567 10471 4573
rect 10594 4564 10600 4576
rect 10652 4564 10658 4616
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9769 4471 9827 4477
rect 9769 4468 9781 4471
rect 9732 4440 9781 4468
rect 9732 4428 9738 4440
rect 9769 4437 9781 4440
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 10505 4471 10563 4477
rect 10505 4437 10517 4471
rect 10551 4468 10563 4471
rect 10686 4468 10692 4480
rect 10551 4440 10692 4468
rect 10551 4437 10563 4440
rect 10505 4431 10563 4437
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11532 4468 11560 4644
rect 11716 4644 12204 4672
rect 12268 4644 12357 4672
rect 11716 4613 11744 4644
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 12176 4604 12204 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12452 4644 13124 4672
rect 12452 4604 12480 4644
rect 12176 4576 12480 4604
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 12526 4536 12532 4548
rect 12023 4508 12532 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 12526 4496 12532 4508
rect 12584 4496 12590 4548
rect 13096 4536 13124 4644
rect 13464 4613 13492 4712
rect 13556 4681 13584 4780
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15105 4811 15163 4817
rect 15105 4808 15117 4811
rect 14976 4780 15117 4808
rect 14976 4768 14982 4780
rect 15105 4777 15117 4780
rect 15151 4808 15163 4811
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 15151 4780 17785 4808
rect 15151 4777 15163 4780
rect 15105 4771 15163 4777
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 27430 4808 27436 4820
rect 17773 4771 17831 4777
rect 26068 4780 27436 4808
rect 13814 4700 13820 4752
rect 13872 4700 13878 4752
rect 15930 4700 15936 4752
rect 15988 4740 15994 4752
rect 15988 4712 16528 4740
rect 15988 4700 15994 4712
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4641 13599 4675
rect 13541 4635 13599 4641
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4641 13783 4675
rect 13832 4672 13860 4700
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 13832 4644 14289 4672
rect 13725 4635 13783 4641
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 14277 4635 14335 4641
rect 13449 4607 13507 4613
rect 13449 4573 13461 4607
rect 13495 4573 13507 4607
rect 13740 4604 13768 4635
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16080 4644 16436 4672
rect 16080 4632 16086 4644
rect 14182 4604 14188 4616
rect 13740 4576 14188 4604
rect 13449 4567 13507 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 14424 4576 15025 4604
rect 14424 4564 14430 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15286 4564 15292 4616
rect 15344 4564 15350 4616
rect 16408 4613 16436 4644
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 16393 4607 16451 4613
rect 15795 4576 16068 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 15488 4536 15516 4567
rect 13096 4508 15516 4536
rect 12894 4468 12900 4480
rect 11532 4440 12900 4468
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 12986 4428 12992 4480
rect 13044 4428 13050 4480
rect 14918 4428 14924 4480
rect 14976 4428 14982 4480
rect 15930 4428 15936 4480
rect 15988 4428 15994 4480
rect 16040 4477 16068 4576
rect 16393 4573 16405 4607
rect 16439 4573 16451 4607
rect 16393 4567 16451 4573
rect 16500 4536 16528 4712
rect 16574 4632 16580 4684
rect 16632 4632 16638 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17052 4644 18153 4672
rect 17052 4613 17080 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 17402 4564 17408 4616
rect 17460 4564 17466 4616
rect 17678 4564 17684 4616
rect 17736 4564 17742 4616
rect 17770 4564 17776 4616
rect 17828 4604 17834 4616
rect 26068 4613 26096 4780
rect 27430 4768 27436 4780
rect 27488 4768 27494 4820
rect 26605 4743 26663 4749
rect 26605 4709 26617 4743
rect 26651 4740 26663 4743
rect 26651 4712 27016 4740
rect 26651 4709 26663 4712
rect 26605 4703 26663 4709
rect 26988 4681 27016 4712
rect 26973 4675 27031 4681
rect 26973 4641 26985 4675
rect 27019 4641 27031 4675
rect 26973 4635 27031 4641
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17828 4576 17969 4604
rect 17828 4564 17834 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 26053 4607 26111 4613
rect 26053 4573 26065 4607
rect 26099 4573 26111 4607
rect 26053 4567 26111 4573
rect 26234 4564 26240 4616
rect 26292 4564 26298 4616
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4604 26479 4607
rect 27154 4604 27160 4616
rect 26467 4576 27160 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 28353 4607 28411 4613
rect 28353 4573 28365 4607
rect 28399 4604 28411 4607
rect 28718 4604 28724 4616
rect 28399 4576 28724 4604
rect 28399 4573 28411 4576
rect 28353 4567 28411 4573
rect 28718 4564 28724 4576
rect 28776 4564 28782 4616
rect 17221 4539 17279 4545
rect 17221 4536 17233 4539
rect 16500 4508 17233 4536
rect 17221 4505 17233 4508
rect 17267 4505 17279 4539
rect 17221 4499 17279 4505
rect 17313 4539 17371 4545
rect 17313 4505 17325 4539
rect 17359 4536 17371 4539
rect 18414 4536 18420 4548
rect 17359 4508 18420 4536
rect 17359 4505 17371 4508
rect 17313 4499 17371 4505
rect 18414 4496 18420 4508
rect 18472 4496 18478 4548
rect 26329 4539 26387 4545
rect 26329 4505 26341 4539
rect 26375 4536 26387 4539
rect 27709 4539 27767 4545
rect 27709 4536 27721 4539
rect 26375 4508 27721 4536
rect 26375 4505 26387 4508
rect 26329 4499 26387 4505
rect 27709 4505 27721 4508
rect 27755 4505 27767 4539
rect 27709 4499 27767 4505
rect 16025 4471 16083 4477
rect 16025 4437 16037 4471
rect 16071 4437 16083 4471
rect 16025 4431 16083 4437
rect 16485 4471 16543 4477
rect 16485 4437 16497 4471
rect 16531 4468 16543 4471
rect 16666 4468 16672 4480
rect 16531 4440 16672 4468
rect 16531 4437 16543 4440
rect 16485 4431 16543 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17589 4471 17647 4477
rect 17589 4437 17601 4471
rect 17635 4468 17647 4471
rect 17954 4468 17960 4480
rect 17635 4440 17960 4468
rect 17635 4437 17647 4440
rect 17589 4431 17647 4437
rect 17954 4428 17960 4440
rect 18012 4428 18018 4480
rect 27614 4428 27620 4480
rect 27672 4428 27678 4480
rect 1104 4378 31280 4400
rect 1104 4326 4922 4378
rect 4974 4326 4986 4378
rect 5038 4326 5050 4378
rect 5102 4326 5114 4378
rect 5166 4326 5178 4378
rect 5230 4326 5242 4378
rect 5294 4326 10922 4378
rect 10974 4326 10986 4378
rect 11038 4326 11050 4378
rect 11102 4326 11114 4378
rect 11166 4326 11178 4378
rect 11230 4326 11242 4378
rect 11294 4326 16922 4378
rect 16974 4326 16986 4378
rect 17038 4326 17050 4378
rect 17102 4326 17114 4378
rect 17166 4326 17178 4378
rect 17230 4326 17242 4378
rect 17294 4326 22922 4378
rect 22974 4326 22986 4378
rect 23038 4326 23050 4378
rect 23102 4326 23114 4378
rect 23166 4326 23178 4378
rect 23230 4326 23242 4378
rect 23294 4326 28922 4378
rect 28974 4326 28986 4378
rect 29038 4326 29050 4378
rect 29102 4326 29114 4378
rect 29166 4326 29178 4378
rect 29230 4326 29242 4378
rect 29294 4326 31280 4378
rect 1104 4304 31280 4326
rect 15289 4267 15347 4273
rect 15289 4264 15301 4267
rect 14568 4236 15301 4264
rect 14568 4196 14596 4236
rect 15289 4233 15301 4236
rect 15335 4233 15347 4267
rect 15289 4227 15347 4233
rect 16666 4224 16672 4276
rect 16724 4264 16730 4276
rect 16853 4267 16911 4273
rect 16853 4264 16865 4267
rect 16724 4236 16865 4264
rect 16724 4224 16730 4236
rect 16853 4233 16865 4236
rect 16899 4233 16911 4267
rect 16853 4227 16911 4233
rect 18414 4224 18420 4276
rect 18472 4224 18478 4276
rect 9324 4168 9720 4196
rect 14398 4168 14596 4196
rect 14829 4199 14887 4205
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9324 4137 9352 4168
rect 9582 4137 9588 4140
rect 9309 4131 9367 4137
rect 9309 4128 9321 4131
rect 9272 4100 9321 4128
rect 9272 4088 9278 4100
rect 9309 4097 9321 4100
rect 9355 4097 9367 4131
rect 9576 4128 9588 4137
rect 9543 4100 9588 4128
rect 9309 4091 9367 4097
rect 9576 4091 9588 4100
rect 9582 4088 9588 4091
rect 9640 4088 9646 4140
rect 9692 4128 9720 4168
rect 14829 4165 14841 4199
rect 14875 4196 14887 4199
rect 14918 4196 14924 4208
rect 14875 4168 14924 4196
rect 14875 4165 14887 4168
rect 14829 4159 14887 4165
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 27706 4156 27712 4208
rect 27764 4156 27770 4208
rect 11882 4128 11888 4140
rect 9692 4100 11888 4128
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 12152 4131 12210 4137
rect 12152 4097 12164 4131
rect 12198 4128 12210 4131
rect 12434 4128 12440 4140
rect 12198 4100 12440 4128
rect 12198 4097 12210 4100
rect 12152 4091 12210 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 13814 4088 13820 4140
rect 13872 4088 13878 4140
rect 15105 4131 15163 4137
rect 15105 4097 15117 4131
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 13832 4060 13860 4088
rect 13412 4032 13860 4060
rect 13412 4020 13418 4032
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 15120 4060 15148 4091
rect 14884 4032 15148 4060
rect 14884 4020 14890 4032
rect 10689 3995 10747 4001
rect 10689 3961 10701 3995
rect 10735 3992 10747 3995
rect 11422 3992 11428 4004
rect 10735 3964 11428 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 15396 3936 15424 4091
rect 17126 4088 17132 4140
rect 17184 4128 17190 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 17184 4100 17509 4128
rect 17184 4088 17190 4100
rect 17497 4097 17509 4100
rect 17543 4128 17555 4131
rect 17678 4128 17684 4140
rect 17543 4100 17684 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 18233 4131 18291 4137
rect 18233 4128 18245 4131
rect 18012 4100 18245 4128
rect 18012 4088 18018 4100
rect 18233 4097 18245 4100
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 25556 4100 26985 4128
rect 25556 4088 25562 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 19061 4063 19119 4069
rect 19061 4029 19073 4063
rect 19107 4060 19119 4063
rect 19426 4060 19432 4072
rect 19107 4032 19432 4060
rect 19107 4029 19119 4032
rect 19061 4023 19119 4029
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 27249 4063 27307 4069
rect 27249 4029 27261 4063
rect 27295 4060 27307 4063
rect 27614 4060 27620 4072
rect 27295 4032 27620 4060
rect 27295 4029 27307 4032
rect 27249 4023 27307 4029
rect 27614 4020 27620 4032
rect 27672 4020 27678 4072
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 14366 3924 14372 3936
rect 13311 3896 14372 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 15378 3884 15384 3936
rect 15436 3884 15442 3936
rect 17678 3884 17684 3936
rect 17736 3884 17742 3936
rect 28718 3884 28724 3936
rect 28776 3884 28782 3936
rect 1104 3834 31280 3856
rect 1104 3782 4182 3834
rect 4234 3782 4246 3834
rect 4298 3782 4310 3834
rect 4362 3782 4374 3834
rect 4426 3782 4438 3834
rect 4490 3782 4502 3834
rect 4554 3782 10182 3834
rect 10234 3782 10246 3834
rect 10298 3782 10310 3834
rect 10362 3782 10374 3834
rect 10426 3782 10438 3834
rect 10490 3782 10502 3834
rect 10554 3782 16182 3834
rect 16234 3782 16246 3834
rect 16298 3782 16310 3834
rect 16362 3782 16374 3834
rect 16426 3782 16438 3834
rect 16490 3782 16502 3834
rect 16554 3782 22182 3834
rect 22234 3782 22246 3834
rect 22298 3782 22310 3834
rect 22362 3782 22374 3834
rect 22426 3782 22438 3834
rect 22490 3782 22502 3834
rect 22554 3782 28182 3834
rect 28234 3782 28246 3834
rect 28298 3782 28310 3834
rect 28362 3782 28374 3834
rect 28426 3782 28438 3834
rect 28490 3782 28502 3834
rect 28554 3782 31280 3834
rect 1104 3760 31280 3782
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10744 3692 10885 3720
rect 10744 3680 10750 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 12526 3680 12532 3732
rect 12584 3720 12590 3732
rect 14093 3723 14151 3729
rect 14093 3720 14105 3723
rect 12584 3692 14105 3720
rect 12584 3680 12590 3692
rect 14093 3689 14105 3692
rect 14139 3689 14151 3723
rect 14093 3683 14151 3689
rect 15764 3692 16804 3720
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 10827 3624 11560 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 9214 3544 9220 3596
rect 9272 3544 9278 3596
rect 11532 3593 11560 3624
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3584 11575 3587
rect 11698 3584 11704 3596
rect 11563 3556 11704 3584
rect 11563 3553 11575 3556
rect 11517 3547 11575 3553
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 11900 3584 11928 3680
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 11900 3556 12173 3584
rect 12161 3553 12173 3556
rect 12207 3553 12219 3587
rect 12161 3547 12219 3553
rect 12437 3587 12495 3593
rect 12437 3553 12449 3587
rect 12483 3584 12495 3587
rect 12986 3584 12992 3596
rect 12483 3556 12992 3584
rect 12483 3553 12495 3556
rect 12437 3547 12495 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14645 3587 14703 3593
rect 14645 3584 14657 3587
rect 13964 3556 14657 3584
rect 13964 3544 13970 3556
rect 14645 3553 14657 3556
rect 14691 3553 14703 3587
rect 14645 3547 14703 3553
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 15764 3593 15792 3692
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 14884 3556 15761 3584
rect 14884 3544 14890 3556
rect 15749 3553 15761 3556
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 9232 3516 9260 3544
rect 9401 3519 9459 3525
rect 9401 3516 9413 3519
rect 9232 3488 9413 3516
rect 9401 3485 9413 3488
rect 9447 3485 9459 3519
rect 9401 3479 9459 3485
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 16016 3519 16074 3525
rect 16016 3485 16028 3519
rect 16062 3485 16074 3519
rect 16776 3516 16804 3692
rect 17126 3680 17132 3732
rect 17184 3680 17190 3732
rect 27249 3723 27307 3729
rect 27249 3689 27261 3723
rect 27295 3720 27307 3723
rect 27706 3720 27712 3732
rect 27295 3692 27712 3720
rect 27295 3689 27307 3692
rect 27249 3683 27307 3689
rect 27706 3680 27712 3692
rect 27764 3680 27770 3732
rect 27338 3612 27344 3664
rect 27396 3612 27402 3664
rect 17589 3587 17647 3593
rect 17589 3553 17601 3587
rect 17635 3584 17647 3587
rect 17678 3584 17684 3596
rect 17635 3556 17684 3584
rect 17635 3553 17647 3556
rect 17589 3547 17647 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 18708 3556 19349 3584
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 16776 3488 17325 3516
rect 16016 3479 16074 3485
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 18708 3502 18736 3556
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 19337 3547 19395 3553
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 17313 3479 17371 3485
rect 18892 3488 19441 3516
rect 9668 3451 9726 3457
rect 9668 3417 9680 3451
rect 9714 3448 9726 3451
rect 9766 3448 9772 3460
rect 9714 3420 9772 3448
rect 9714 3417 9726 3420
rect 9668 3411 9726 3417
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 14921 3451 14979 3457
rect 14921 3448 14933 3451
rect 13662 3420 14933 3448
rect 14921 3417 14933 3420
rect 14967 3417 14979 3451
rect 14921 3411 14979 3417
rect 15028 3380 15056 3479
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16040 3448 16068 3479
rect 15988 3420 16068 3448
rect 15988 3408 15994 3420
rect 15378 3380 15384 3392
rect 15028 3352 15384 3380
rect 15378 3340 15384 3352
rect 15436 3380 15442 3392
rect 18892 3380 18920 3488
rect 19429 3485 19441 3488
rect 19475 3516 19487 3519
rect 27157 3519 27215 3525
rect 27157 3516 27169 3519
rect 19475 3488 27169 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 27157 3485 27169 3488
rect 27203 3516 27215 3519
rect 27356 3516 27384 3612
rect 27203 3488 27384 3516
rect 27203 3485 27215 3488
rect 27157 3479 27215 3485
rect 15436 3352 18920 3380
rect 19061 3383 19119 3389
rect 15436 3340 15442 3352
rect 19061 3349 19073 3383
rect 19107 3380 19119 3383
rect 19426 3380 19432 3392
rect 19107 3352 19432 3380
rect 19107 3349 19119 3352
rect 19061 3343 19119 3349
rect 19426 3340 19432 3352
rect 19484 3380 19490 3392
rect 20254 3380 20260 3392
rect 19484 3352 20260 3380
rect 19484 3340 19490 3352
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 1104 3290 31280 3312
rect 1104 3238 4922 3290
rect 4974 3238 4986 3290
rect 5038 3238 5050 3290
rect 5102 3238 5114 3290
rect 5166 3238 5178 3290
rect 5230 3238 5242 3290
rect 5294 3238 10922 3290
rect 10974 3238 10986 3290
rect 11038 3238 11050 3290
rect 11102 3238 11114 3290
rect 11166 3238 11178 3290
rect 11230 3238 11242 3290
rect 11294 3238 16922 3290
rect 16974 3238 16986 3290
rect 17038 3238 17050 3290
rect 17102 3238 17114 3290
rect 17166 3238 17178 3290
rect 17230 3238 17242 3290
rect 17294 3238 22922 3290
rect 22974 3238 22986 3290
rect 23038 3238 23050 3290
rect 23102 3238 23114 3290
rect 23166 3238 23178 3290
rect 23230 3238 23242 3290
rect 23294 3238 28922 3290
rect 28974 3238 28986 3290
rect 29038 3238 29050 3290
rect 29102 3238 29114 3290
rect 29166 3238 29178 3290
rect 29230 3238 29242 3290
rect 29294 3238 31280 3290
rect 1104 3216 31280 3238
rect 1104 2746 31280 2768
rect 1104 2694 4182 2746
rect 4234 2694 4246 2746
rect 4298 2694 4310 2746
rect 4362 2694 4374 2746
rect 4426 2694 4438 2746
rect 4490 2694 4502 2746
rect 4554 2694 10182 2746
rect 10234 2694 10246 2746
rect 10298 2694 10310 2746
rect 10362 2694 10374 2746
rect 10426 2694 10438 2746
rect 10490 2694 10502 2746
rect 10554 2694 16182 2746
rect 16234 2694 16246 2746
rect 16298 2694 16310 2746
rect 16362 2694 16374 2746
rect 16426 2694 16438 2746
rect 16490 2694 16502 2746
rect 16554 2694 22182 2746
rect 22234 2694 22246 2746
rect 22298 2694 22310 2746
rect 22362 2694 22374 2746
rect 22426 2694 22438 2746
rect 22490 2694 22502 2746
rect 22554 2694 28182 2746
rect 28234 2694 28246 2746
rect 28298 2694 28310 2746
rect 28362 2694 28374 2746
rect 28426 2694 28438 2746
rect 28490 2694 28502 2746
rect 28554 2694 31280 2746
rect 1104 2672 31280 2694
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 28629 2635 28687 2641
rect 28629 2632 28641 2635
rect 9916 2604 28641 2632
rect 9916 2592 9922 2604
rect 28629 2601 28641 2604
rect 28675 2601 28687 2635
rect 28629 2595 28687 2601
rect 13354 2496 13360 2508
rect 1780 2468 13360 2496
rect 1780 2437 1808 2468
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 13906 2428 13912 2440
rect 5491 2400 13912 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2428 17095 2431
rect 19150 2428 19156 2440
rect 17083 2400 19156 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 20254 2388 20260 2440
rect 20312 2428 20318 2440
rect 22741 2431 22799 2437
rect 22741 2428 22753 2431
rect 20312 2400 22753 2428
rect 20312 2388 20318 2400
rect 22741 2397 22753 2400
rect 22787 2397 22799 2431
rect 22741 2391 22799 2397
rect 28718 2388 28724 2440
rect 28776 2428 28782 2440
rect 30653 2431 30711 2437
rect 30653 2428 30665 2431
rect 28776 2400 30665 2428
rect 28776 2388 28782 2400
rect 30653 2397 30665 2400
rect 30699 2397 30711 2431
rect 30653 2391 30711 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 10870 2320 10876 2372
rect 10928 2320 10934 2372
rect 11241 2363 11299 2369
rect 11241 2329 11253 2363
rect 11287 2360 11299 2363
rect 13262 2360 13268 2372
rect 11287 2332 13268 2360
rect 11287 2329 11299 2332
rect 11241 2323 11299 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 28534 2320 28540 2372
rect 28592 2320 28598 2372
rect 5350 2252 5356 2304
rect 5408 2252 5414 2304
rect 16758 2252 16764 2304
rect 16816 2252 16822 2304
rect 22554 2252 22560 2304
rect 22612 2292 22618 2304
rect 22833 2295 22891 2301
rect 22833 2292 22845 2295
rect 22612 2264 22845 2292
rect 22612 2252 22618 2264
rect 22833 2261 22845 2264
rect 22879 2261 22891 2295
rect 22833 2255 22891 2261
rect 30834 2252 30840 2304
rect 30892 2252 30898 2304
rect 1104 2202 31280 2224
rect 1104 2150 4922 2202
rect 4974 2150 4986 2202
rect 5038 2150 5050 2202
rect 5102 2150 5114 2202
rect 5166 2150 5178 2202
rect 5230 2150 5242 2202
rect 5294 2150 10922 2202
rect 10974 2150 10986 2202
rect 11038 2150 11050 2202
rect 11102 2150 11114 2202
rect 11166 2150 11178 2202
rect 11230 2150 11242 2202
rect 11294 2150 16922 2202
rect 16974 2150 16986 2202
rect 17038 2150 17050 2202
rect 17102 2150 17114 2202
rect 17166 2150 17178 2202
rect 17230 2150 17242 2202
rect 17294 2150 22922 2202
rect 22974 2150 22986 2202
rect 23038 2150 23050 2202
rect 23102 2150 23114 2202
rect 23166 2150 23178 2202
rect 23230 2150 23242 2202
rect 23294 2150 28922 2202
rect 28974 2150 28986 2202
rect 29038 2150 29050 2202
rect 29102 2150 29114 2202
rect 29166 2150 29178 2202
rect 29230 2150 29242 2202
rect 29294 2150 31280 2202
rect 1104 2128 31280 2150
<< via1 >>
rect 4182 32070 4234 32122
rect 4246 32070 4298 32122
rect 4310 32070 4362 32122
rect 4374 32070 4426 32122
rect 4438 32070 4490 32122
rect 4502 32070 4554 32122
rect 10182 32070 10234 32122
rect 10246 32070 10298 32122
rect 10310 32070 10362 32122
rect 10374 32070 10426 32122
rect 10438 32070 10490 32122
rect 10502 32070 10554 32122
rect 16182 32070 16234 32122
rect 16246 32070 16298 32122
rect 16310 32070 16362 32122
rect 16374 32070 16426 32122
rect 16438 32070 16490 32122
rect 16502 32070 16554 32122
rect 22182 32070 22234 32122
rect 22246 32070 22298 32122
rect 22310 32070 22362 32122
rect 22374 32070 22426 32122
rect 22438 32070 22490 32122
rect 22502 32070 22554 32122
rect 28182 32070 28234 32122
rect 28246 32070 28298 32122
rect 28310 32070 28362 32122
rect 28374 32070 28426 32122
rect 28438 32070 28490 32122
rect 28502 32070 28554 32122
rect 18052 31968 18104 32020
rect 23848 31968 23900 32020
rect 18788 31900 18840 31952
rect 1308 31764 1360 31816
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 7104 31764 7156 31816
rect 12256 31764 12308 31816
rect 18144 31807 18196 31816
rect 18144 31773 18153 31807
rect 18153 31773 18187 31807
rect 18187 31773 18196 31807
rect 18144 31764 18196 31773
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 24492 31807 24544 31816
rect 24492 31773 24501 31807
rect 24501 31773 24535 31807
rect 24535 31773 24544 31807
rect 24492 31764 24544 31773
rect 29644 31764 29696 31816
rect 12532 31671 12584 31680
rect 12532 31637 12541 31671
rect 12541 31637 12575 31671
rect 12575 31637 12584 31671
rect 12532 31628 12584 31637
rect 18328 31671 18380 31680
rect 18328 31637 18337 31671
rect 18337 31637 18371 31671
rect 18371 31637 18380 31671
rect 18328 31628 18380 31637
rect 26700 31628 26752 31680
rect 4922 31526 4974 31578
rect 4986 31526 5038 31578
rect 5050 31526 5102 31578
rect 5114 31526 5166 31578
rect 5178 31526 5230 31578
rect 5242 31526 5294 31578
rect 10922 31526 10974 31578
rect 10986 31526 11038 31578
rect 11050 31526 11102 31578
rect 11114 31526 11166 31578
rect 11178 31526 11230 31578
rect 11242 31526 11294 31578
rect 16922 31526 16974 31578
rect 16986 31526 17038 31578
rect 17050 31526 17102 31578
rect 17114 31526 17166 31578
rect 17178 31526 17230 31578
rect 17242 31526 17294 31578
rect 22922 31526 22974 31578
rect 22986 31526 23038 31578
rect 23050 31526 23102 31578
rect 23114 31526 23166 31578
rect 23178 31526 23230 31578
rect 23242 31526 23294 31578
rect 28922 31526 28974 31578
rect 28986 31526 29038 31578
rect 29050 31526 29102 31578
rect 29114 31526 29166 31578
rect 29178 31526 29230 31578
rect 29242 31526 29294 31578
rect 18328 31424 18380 31476
rect 8576 31220 8628 31272
rect 9128 31220 9180 31272
rect 12532 31356 12584 31408
rect 21088 31356 21140 31408
rect 20720 31331 20772 31340
rect 20720 31297 20729 31331
rect 20729 31297 20763 31331
rect 20763 31297 20772 31331
rect 20720 31288 20772 31297
rect 21364 31331 21416 31340
rect 21364 31297 21373 31331
rect 21373 31297 21407 31331
rect 21407 31297 21416 31331
rect 21364 31288 21416 31297
rect 24216 31288 24268 31340
rect 12900 31263 12952 31272
rect 12900 31229 12909 31263
rect 12909 31229 12943 31263
rect 12943 31229 12952 31263
rect 12900 31220 12952 31229
rect 17960 31220 18012 31272
rect 14556 31152 14608 31204
rect 16948 31152 17000 31204
rect 18696 31220 18748 31272
rect 19800 31263 19852 31272
rect 19800 31229 19809 31263
rect 19809 31229 19843 31263
rect 19843 31229 19852 31263
rect 19800 31220 19852 31229
rect 21640 31220 21692 31272
rect 23296 31263 23348 31272
rect 23296 31229 23305 31263
rect 23305 31229 23339 31263
rect 23339 31229 23348 31263
rect 23296 31220 23348 31229
rect 24676 31263 24728 31272
rect 24676 31229 24685 31263
rect 24685 31229 24719 31263
rect 24719 31229 24728 31263
rect 24676 31220 24728 31229
rect 7012 31127 7064 31136
rect 7012 31093 7021 31127
rect 7021 31093 7055 31127
rect 7055 31093 7064 31127
rect 7012 31084 7064 31093
rect 10968 31127 11020 31136
rect 10968 31093 10977 31127
rect 10977 31093 11011 31127
rect 11011 31093 11020 31127
rect 10968 31084 11020 31093
rect 17592 31127 17644 31136
rect 17592 31093 17601 31127
rect 17601 31093 17635 31127
rect 17635 31093 17644 31127
rect 17592 31084 17644 31093
rect 20536 31127 20588 31136
rect 20536 31093 20545 31127
rect 20545 31093 20579 31127
rect 20579 31093 20588 31127
rect 20536 31084 20588 31093
rect 21548 31127 21600 31136
rect 21548 31093 21557 31127
rect 21557 31093 21591 31127
rect 21591 31093 21600 31127
rect 21548 31084 21600 31093
rect 21824 31127 21876 31136
rect 21824 31093 21833 31127
rect 21833 31093 21867 31127
rect 21867 31093 21876 31127
rect 21824 31084 21876 31093
rect 22744 31127 22796 31136
rect 22744 31093 22753 31127
rect 22753 31093 22787 31127
rect 22787 31093 22796 31127
rect 22744 31084 22796 31093
rect 24032 31127 24084 31136
rect 24032 31093 24041 31127
rect 24041 31093 24075 31127
rect 24075 31093 24084 31127
rect 24032 31084 24084 31093
rect 24124 31127 24176 31136
rect 24124 31093 24133 31127
rect 24133 31093 24167 31127
rect 24167 31093 24176 31127
rect 24124 31084 24176 31093
rect 4182 30982 4234 31034
rect 4246 30982 4298 31034
rect 4310 30982 4362 31034
rect 4374 30982 4426 31034
rect 4438 30982 4490 31034
rect 4502 30982 4554 31034
rect 10182 30982 10234 31034
rect 10246 30982 10298 31034
rect 10310 30982 10362 31034
rect 10374 30982 10426 31034
rect 10438 30982 10490 31034
rect 10502 30982 10554 31034
rect 16182 30982 16234 31034
rect 16246 30982 16298 31034
rect 16310 30982 16362 31034
rect 16374 30982 16426 31034
rect 16438 30982 16490 31034
rect 16502 30982 16554 31034
rect 22182 30982 22234 31034
rect 22246 30982 22298 31034
rect 22310 30982 22362 31034
rect 22374 30982 22426 31034
rect 22438 30982 22490 31034
rect 22502 30982 22554 31034
rect 28182 30982 28234 31034
rect 28246 30982 28298 31034
rect 28310 30982 28362 31034
rect 28374 30982 28426 31034
rect 28438 30982 28490 31034
rect 28502 30982 28554 31034
rect 12900 30880 12952 30932
rect 16948 30880 17000 30932
rect 10416 30812 10468 30864
rect 9680 30744 9732 30796
rect 5632 30676 5684 30728
rect 7380 30719 7432 30728
rect 7380 30685 7389 30719
rect 7389 30685 7423 30719
rect 7423 30685 7432 30719
rect 7380 30676 7432 30685
rect 8116 30608 8168 30660
rect 8576 30540 8628 30592
rect 10048 30676 10100 30728
rect 10968 30719 11020 30728
rect 10968 30685 11002 30719
rect 11002 30685 11020 30719
rect 10968 30676 11020 30685
rect 14004 30676 14056 30728
rect 14648 30676 14700 30728
rect 11888 30608 11940 30660
rect 12808 30608 12860 30660
rect 8944 30583 8996 30592
rect 8944 30549 8953 30583
rect 8953 30549 8987 30583
rect 8987 30549 8996 30583
rect 8944 30540 8996 30549
rect 9128 30540 9180 30592
rect 12072 30540 12124 30592
rect 12348 30540 12400 30592
rect 15016 30540 15068 30592
rect 17592 30880 17644 30932
rect 19800 30880 19852 30932
rect 21548 30880 21600 30932
rect 22836 30880 22888 30932
rect 23296 30880 23348 30932
rect 24124 30880 24176 30932
rect 24216 30923 24268 30932
rect 24216 30889 24225 30923
rect 24225 30889 24259 30923
rect 24259 30889 24268 30923
rect 24216 30880 24268 30889
rect 24676 30880 24728 30932
rect 17316 30719 17368 30728
rect 17316 30685 17325 30719
rect 17325 30685 17359 30719
rect 17359 30685 17368 30719
rect 17316 30676 17368 30685
rect 19984 30676 20036 30728
rect 24952 30676 25004 30728
rect 15568 30583 15620 30592
rect 15568 30549 15577 30583
rect 15577 30549 15611 30583
rect 15611 30549 15620 30583
rect 15568 30540 15620 30549
rect 20536 30651 20588 30660
rect 20536 30617 20570 30651
rect 20570 30617 20588 30651
rect 20536 30608 20588 30617
rect 21088 30608 21140 30660
rect 17408 30540 17460 30592
rect 21640 30583 21692 30592
rect 21640 30549 21649 30583
rect 21649 30549 21683 30583
rect 21683 30549 21692 30583
rect 21640 30540 21692 30549
rect 23664 30608 23716 30660
rect 24032 30608 24084 30660
rect 26700 30540 26752 30592
rect 4922 30438 4974 30490
rect 4986 30438 5038 30490
rect 5050 30438 5102 30490
rect 5114 30438 5166 30490
rect 5178 30438 5230 30490
rect 5242 30438 5294 30490
rect 10922 30438 10974 30490
rect 10986 30438 11038 30490
rect 11050 30438 11102 30490
rect 11114 30438 11166 30490
rect 11178 30438 11230 30490
rect 11242 30438 11294 30490
rect 16922 30438 16974 30490
rect 16986 30438 17038 30490
rect 17050 30438 17102 30490
rect 17114 30438 17166 30490
rect 17178 30438 17230 30490
rect 17242 30438 17294 30490
rect 22922 30438 22974 30490
rect 22986 30438 23038 30490
rect 23050 30438 23102 30490
rect 23114 30438 23166 30490
rect 23178 30438 23230 30490
rect 23242 30438 23294 30490
rect 28922 30438 28974 30490
rect 28986 30438 29038 30490
rect 29050 30438 29102 30490
rect 29114 30438 29166 30490
rect 29178 30438 29230 30490
rect 29242 30438 29294 30490
rect 5632 30336 5684 30388
rect 7012 30336 7064 30388
rect 8116 30379 8168 30388
rect 8116 30345 8125 30379
rect 8125 30345 8159 30379
rect 8159 30345 8168 30379
rect 8116 30336 8168 30345
rect 8944 30336 8996 30388
rect 940 30200 992 30252
rect 8024 30200 8076 30252
rect 11888 30311 11940 30320
rect 11888 30277 11897 30311
rect 11897 30277 11931 30311
rect 11931 30277 11940 30311
rect 11888 30268 11940 30277
rect 12256 30336 12308 30388
rect 14004 30379 14056 30388
rect 14004 30345 14013 30379
rect 14013 30345 14047 30379
rect 14047 30345 14056 30379
rect 14004 30336 14056 30345
rect 15568 30336 15620 30388
rect 17408 30336 17460 30388
rect 18696 30336 18748 30388
rect 11520 30200 11572 30252
rect 6000 30064 6052 30116
rect 10416 30132 10468 30184
rect 10784 30132 10836 30184
rect 12348 30243 12400 30252
rect 12348 30209 12357 30243
rect 12357 30209 12391 30243
rect 12391 30209 12400 30243
rect 12348 30200 12400 30209
rect 17316 30200 17368 30252
rect 14556 30175 14608 30184
rect 14556 30141 14565 30175
rect 14565 30141 14599 30175
rect 14599 30141 14608 30175
rect 14556 30132 14608 30141
rect 20720 30336 20772 30388
rect 21824 30336 21876 30388
rect 22744 30336 22796 30388
rect 19984 30268 20036 30320
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 22100 30200 22152 30252
rect 23020 30243 23072 30252
rect 23020 30209 23029 30243
rect 23029 30209 23063 30243
rect 23063 30209 23072 30243
rect 23020 30200 23072 30209
rect 23204 30200 23256 30252
rect 24952 30268 25004 30320
rect 11520 30107 11572 30116
rect 11520 30073 11529 30107
rect 11529 30073 11563 30107
rect 11563 30073 11572 30107
rect 11520 30064 11572 30073
rect 12808 29996 12860 30048
rect 18880 30064 18932 30116
rect 17960 29996 18012 30048
rect 20904 29996 20956 30048
rect 21364 29996 21416 30048
rect 23112 29996 23164 30048
rect 24768 30039 24820 30048
rect 24768 30005 24777 30039
rect 24777 30005 24811 30039
rect 24811 30005 24820 30039
rect 24768 29996 24820 30005
rect 4182 29894 4234 29946
rect 4246 29894 4298 29946
rect 4310 29894 4362 29946
rect 4374 29894 4426 29946
rect 4438 29894 4490 29946
rect 4502 29894 4554 29946
rect 10182 29894 10234 29946
rect 10246 29894 10298 29946
rect 10310 29894 10362 29946
rect 10374 29894 10426 29946
rect 10438 29894 10490 29946
rect 10502 29894 10554 29946
rect 16182 29894 16234 29946
rect 16246 29894 16298 29946
rect 16310 29894 16362 29946
rect 16374 29894 16426 29946
rect 16438 29894 16490 29946
rect 16502 29894 16554 29946
rect 22182 29894 22234 29946
rect 22246 29894 22298 29946
rect 22310 29894 22362 29946
rect 22374 29894 22426 29946
rect 22438 29894 22490 29946
rect 22502 29894 22554 29946
rect 28182 29894 28234 29946
rect 28246 29894 28298 29946
rect 28310 29894 28362 29946
rect 28374 29894 28426 29946
rect 28438 29894 28490 29946
rect 28502 29894 28554 29946
rect 11980 29792 12032 29844
rect 15292 29792 15344 29844
rect 23020 29792 23072 29844
rect 24768 29792 24820 29844
rect 21916 29724 21968 29776
rect 8484 29631 8536 29640
rect 8484 29597 8493 29631
rect 8493 29597 8527 29631
rect 8527 29597 8536 29631
rect 8484 29588 8536 29597
rect 10048 29588 10100 29640
rect 11336 29588 11388 29640
rect 12348 29631 12400 29640
rect 12348 29597 12357 29631
rect 12357 29597 12391 29631
rect 12391 29597 12400 29631
rect 12348 29588 12400 29597
rect 14648 29631 14700 29640
rect 14648 29597 14657 29631
rect 14657 29597 14691 29631
rect 14691 29597 14700 29631
rect 14648 29588 14700 29597
rect 12256 29520 12308 29572
rect 14924 29563 14976 29572
rect 14924 29529 14958 29563
rect 14958 29529 14976 29563
rect 14924 29520 14976 29529
rect 8300 29495 8352 29504
rect 8300 29461 8309 29495
rect 8309 29461 8343 29495
rect 8343 29461 8352 29495
rect 8300 29452 8352 29461
rect 9312 29452 9364 29504
rect 9404 29495 9456 29504
rect 9404 29461 9413 29495
rect 9413 29461 9447 29495
rect 9447 29461 9456 29495
rect 9404 29452 9456 29461
rect 10692 29495 10744 29504
rect 10692 29461 10701 29495
rect 10701 29461 10735 29495
rect 10735 29461 10744 29495
rect 10692 29452 10744 29461
rect 11704 29495 11756 29504
rect 11704 29461 11713 29495
rect 11713 29461 11747 29495
rect 11747 29461 11756 29495
rect 11704 29452 11756 29461
rect 12532 29452 12584 29504
rect 15384 29520 15436 29572
rect 16028 29588 16080 29640
rect 17316 29588 17368 29640
rect 18880 29588 18932 29640
rect 19340 29520 19392 29572
rect 19892 29588 19944 29640
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 23940 29724 23992 29776
rect 24400 29724 24452 29776
rect 24492 29656 24544 29708
rect 23112 29631 23164 29640
rect 23112 29597 23121 29631
rect 23121 29597 23155 29631
rect 23155 29597 23164 29631
rect 23112 29588 23164 29597
rect 24952 29656 25004 29708
rect 19616 29563 19668 29572
rect 19616 29529 19625 29563
rect 19625 29529 19659 29563
rect 19659 29529 19668 29563
rect 19616 29520 19668 29529
rect 26240 29520 26292 29572
rect 15200 29452 15252 29504
rect 16028 29495 16080 29504
rect 16028 29461 16037 29495
rect 16037 29461 16071 29495
rect 16071 29461 16080 29495
rect 16028 29452 16080 29461
rect 16120 29495 16172 29504
rect 16120 29461 16129 29495
rect 16129 29461 16163 29495
rect 16163 29461 16172 29495
rect 16120 29452 16172 29461
rect 20812 29495 20864 29504
rect 20812 29461 20821 29495
rect 20821 29461 20855 29495
rect 20855 29461 20864 29495
rect 20812 29452 20864 29461
rect 23388 29495 23440 29504
rect 23388 29461 23397 29495
rect 23397 29461 23431 29495
rect 23431 29461 23440 29495
rect 23388 29452 23440 29461
rect 23848 29452 23900 29504
rect 24308 29452 24360 29504
rect 24584 29495 24636 29504
rect 24584 29461 24593 29495
rect 24593 29461 24627 29495
rect 24627 29461 24636 29495
rect 24584 29452 24636 29461
rect 4922 29350 4974 29402
rect 4986 29350 5038 29402
rect 5050 29350 5102 29402
rect 5114 29350 5166 29402
rect 5178 29350 5230 29402
rect 5242 29350 5294 29402
rect 10922 29350 10974 29402
rect 10986 29350 11038 29402
rect 11050 29350 11102 29402
rect 11114 29350 11166 29402
rect 11178 29350 11230 29402
rect 11242 29350 11294 29402
rect 16922 29350 16974 29402
rect 16986 29350 17038 29402
rect 17050 29350 17102 29402
rect 17114 29350 17166 29402
rect 17178 29350 17230 29402
rect 17242 29350 17294 29402
rect 22922 29350 22974 29402
rect 22986 29350 23038 29402
rect 23050 29350 23102 29402
rect 23114 29350 23166 29402
rect 23178 29350 23230 29402
rect 23242 29350 23294 29402
rect 28922 29350 28974 29402
rect 28986 29350 29038 29402
rect 29050 29350 29102 29402
rect 29114 29350 29166 29402
rect 29178 29350 29230 29402
rect 29242 29350 29294 29402
rect 8300 29248 8352 29300
rect 9312 29291 9364 29300
rect 9312 29257 9321 29291
rect 9321 29257 9355 29291
rect 9355 29257 9364 29291
rect 9312 29248 9364 29257
rect 11704 29248 11756 29300
rect 12532 29248 12584 29300
rect 14464 29291 14516 29300
rect 7012 29112 7064 29164
rect 7380 29112 7432 29164
rect 10600 29112 10652 29164
rect 14464 29257 14473 29291
rect 14473 29257 14507 29291
rect 14507 29257 14516 29291
rect 14464 29248 14516 29257
rect 14648 29248 14700 29300
rect 14924 29248 14976 29300
rect 6092 29087 6144 29096
rect 6092 29053 6101 29087
rect 6101 29053 6135 29087
rect 6135 29053 6144 29087
rect 6092 29044 6144 29053
rect 9680 29044 9732 29096
rect 11980 29087 12032 29096
rect 11980 29053 11989 29087
rect 11989 29053 12023 29087
rect 12023 29053 12032 29087
rect 11980 29044 12032 29053
rect 12164 29087 12216 29096
rect 12164 29053 12173 29087
rect 12173 29053 12207 29087
rect 12207 29053 12216 29087
rect 12164 29044 12216 29053
rect 12348 29044 12400 29096
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 12900 29112 12952 29121
rect 13176 29112 13228 29164
rect 15292 29248 15344 29300
rect 16120 29248 16172 29300
rect 19432 29180 19484 29232
rect 19800 29248 19852 29300
rect 20720 29248 20772 29300
rect 20812 29248 20864 29300
rect 24584 29248 24636 29300
rect 26240 29291 26292 29300
rect 26240 29257 26249 29291
rect 26249 29257 26283 29291
rect 26283 29257 26292 29291
rect 26240 29248 26292 29257
rect 19616 29180 19668 29232
rect 19800 29155 19852 29164
rect 19800 29121 19809 29155
rect 19809 29121 19843 29155
rect 19843 29121 19852 29155
rect 19800 29112 19852 29121
rect 19892 29155 19944 29164
rect 19892 29121 19901 29155
rect 19901 29121 19935 29155
rect 19935 29121 19944 29155
rect 19892 29112 19944 29121
rect 20352 29112 20404 29164
rect 18880 29044 18932 29096
rect 19340 29087 19392 29096
rect 19340 29053 19349 29087
rect 19349 29053 19383 29087
rect 19383 29053 19392 29087
rect 19340 29044 19392 29053
rect 19984 29044 20036 29096
rect 22836 29044 22888 29096
rect 24400 29155 24452 29164
rect 24400 29121 24409 29155
rect 24409 29121 24443 29155
rect 24443 29121 24452 29155
rect 24400 29112 24452 29121
rect 24676 29112 24728 29164
rect 24492 29044 24544 29096
rect 24952 29087 25004 29096
rect 24952 29053 24961 29087
rect 24961 29053 24995 29087
rect 24995 29053 25004 29087
rect 24952 29044 25004 29053
rect 24308 28976 24360 29028
rect 24676 28976 24728 29028
rect 5540 28951 5592 28960
rect 5540 28917 5549 28951
rect 5549 28917 5583 28951
rect 5583 28917 5592 28951
rect 5540 28908 5592 28917
rect 6368 28951 6420 28960
rect 6368 28917 6377 28951
rect 6377 28917 6411 28951
rect 6411 28917 6420 28951
rect 6368 28908 6420 28917
rect 6460 28908 6512 28960
rect 9128 28908 9180 28960
rect 11520 28951 11572 28960
rect 11520 28917 11529 28951
rect 11529 28917 11563 28951
rect 11563 28917 11572 28951
rect 11520 28908 11572 28917
rect 11612 28908 11664 28960
rect 13084 28908 13136 28960
rect 15108 28908 15160 28960
rect 17684 28951 17736 28960
rect 17684 28917 17693 28951
rect 17693 28917 17727 28951
rect 17727 28917 17736 28951
rect 17684 28908 17736 28917
rect 21824 28951 21876 28960
rect 21824 28917 21833 28951
rect 21833 28917 21867 28951
rect 21867 28917 21876 28951
rect 21824 28908 21876 28917
rect 24032 28951 24084 28960
rect 24032 28917 24041 28951
rect 24041 28917 24075 28951
rect 24075 28917 24084 28951
rect 24032 28908 24084 28917
rect 4182 28806 4234 28858
rect 4246 28806 4298 28858
rect 4310 28806 4362 28858
rect 4374 28806 4426 28858
rect 4438 28806 4490 28858
rect 4502 28806 4554 28858
rect 10182 28806 10234 28858
rect 10246 28806 10298 28858
rect 10310 28806 10362 28858
rect 10374 28806 10426 28858
rect 10438 28806 10490 28858
rect 10502 28806 10554 28858
rect 16182 28806 16234 28858
rect 16246 28806 16298 28858
rect 16310 28806 16362 28858
rect 16374 28806 16426 28858
rect 16438 28806 16490 28858
rect 16502 28806 16554 28858
rect 22182 28806 22234 28858
rect 22246 28806 22298 28858
rect 22310 28806 22362 28858
rect 22374 28806 22426 28858
rect 22438 28806 22490 28858
rect 22502 28806 22554 28858
rect 28182 28806 28234 28858
rect 28246 28806 28298 28858
rect 28310 28806 28362 28858
rect 28374 28806 28426 28858
rect 28438 28806 28490 28858
rect 28502 28806 28554 28858
rect 7012 28747 7064 28756
rect 7012 28713 7021 28747
rect 7021 28713 7055 28747
rect 7055 28713 7064 28747
rect 7012 28704 7064 28713
rect 8484 28704 8536 28756
rect 10600 28704 10652 28756
rect 13176 28704 13228 28756
rect 19800 28704 19852 28756
rect 20996 28704 21048 28756
rect 11336 28636 11388 28688
rect 7380 28568 7432 28620
rect 7472 28568 7524 28620
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 9956 28568 10008 28620
rect 12164 28568 12216 28620
rect 9404 28500 9456 28552
rect 11520 28500 11572 28552
rect 12072 28543 12124 28552
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 12348 28543 12400 28552
rect 12348 28509 12357 28543
rect 12357 28509 12391 28543
rect 12391 28509 12400 28543
rect 12348 28500 12400 28509
rect 6368 28432 6420 28484
rect 8484 28432 8536 28484
rect 11980 28432 12032 28484
rect 12164 28432 12216 28484
rect 13176 28568 13228 28620
rect 14464 28568 14516 28620
rect 8300 28364 8352 28416
rect 15016 28500 15068 28552
rect 15108 28543 15160 28552
rect 15108 28509 15117 28543
rect 15117 28509 15151 28543
rect 15151 28509 15160 28543
rect 15108 28500 15160 28509
rect 15200 28543 15252 28552
rect 15200 28509 15209 28543
rect 15209 28509 15243 28543
rect 15243 28509 15252 28543
rect 15200 28500 15252 28509
rect 15384 28500 15436 28552
rect 15568 28475 15620 28484
rect 15568 28441 15577 28475
rect 15577 28441 15611 28475
rect 15611 28441 15620 28475
rect 15568 28432 15620 28441
rect 15752 28543 15804 28552
rect 15752 28509 15761 28543
rect 15761 28509 15795 28543
rect 15795 28509 15804 28543
rect 15752 28500 15804 28509
rect 17316 28500 17368 28552
rect 18880 28568 18932 28620
rect 20904 28568 20956 28620
rect 20352 28500 20404 28552
rect 21824 28500 21876 28552
rect 17500 28432 17552 28484
rect 14556 28364 14608 28416
rect 15384 28364 15436 28416
rect 19248 28407 19300 28416
rect 19248 28373 19257 28407
rect 19257 28373 19291 28407
rect 19291 28373 19300 28407
rect 19248 28364 19300 28373
rect 19708 28407 19760 28416
rect 19708 28373 19717 28407
rect 19717 28373 19751 28407
rect 19751 28373 19760 28407
rect 19708 28364 19760 28373
rect 22100 28364 22152 28416
rect 4922 28262 4974 28314
rect 4986 28262 5038 28314
rect 5050 28262 5102 28314
rect 5114 28262 5166 28314
rect 5178 28262 5230 28314
rect 5242 28262 5294 28314
rect 10922 28262 10974 28314
rect 10986 28262 11038 28314
rect 11050 28262 11102 28314
rect 11114 28262 11166 28314
rect 11178 28262 11230 28314
rect 11242 28262 11294 28314
rect 16922 28262 16974 28314
rect 16986 28262 17038 28314
rect 17050 28262 17102 28314
rect 17114 28262 17166 28314
rect 17178 28262 17230 28314
rect 17242 28262 17294 28314
rect 22922 28262 22974 28314
rect 22986 28262 23038 28314
rect 23050 28262 23102 28314
rect 23114 28262 23166 28314
rect 23178 28262 23230 28314
rect 23242 28262 23294 28314
rect 28922 28262 28974 28314
rect 28986 28262 29038 28314
rect 29050 28262 29102 28314
rect 29114 28262 29166 28314
rect 29178 28262 29230 28314
rect 29242 28262 29294 28314
rect 5540 28160 5592 28212
rect 6368 28160 6420 28212
rect 6552 28160 6604 28212
rect 8300 28160 8352 28212
rect 8392 28160 8444 28212
rect 15568 28160 15620 28212
rect 17500 28160 17552 28212
rect 4620 28024 4672 28076
rect 13636 28092 13688 28144
rect 6460 28024 6512 28076
rect 7380 28024 7432 28076
rect 7656 28024 7708 28076
rect 6000 27999 6052 28008
rect 6000 27965 6009 27999
rect 6009 27965 6043 27999
rect 6043 27965 6052 27999
rect 6000 27956 6052 27965
rect 8576 28067 8628 28076
rect 8576 28033 8585 28067
rect 8585 28033 8619 28067
rect 8619 28033 8628 28067
rect 8576 28024 8628 28033
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 8760 28024 8812 28033
rect 9128 28024 9180 28076
rect 7748 27931 7800 27940
rect 7748 27897 7757 27931
rect 7757 27897 7791 27931
rect 7791 27897 7800 27931
rect 13728 28024 13780 28076
rect 19248 28160 19300 28212
rect 17684 28092 17736 28144
rect 22284 28092 22336 28144
rect 21640 28024 21692 28076
rect 13544 27956 13596 28008
rect 17316 27956 17368 28008
rect 22468 28024 22520 28076
rect 22652 28024 22704 28076
rect 22928 28067 22980 28076
rect 22928 28033 22937 28067
rect 22937 28033 22971 28067
rect 22971 28033 22980 28067
rect 22928 28024 22980 28033
rect 23388 28024 23440 28076
rect 24032 28024 24084 28076
rect 7748 27888 7800 27897
rect 10692 27888 10744 27940
rect 5356 27863 5408 27872
rect 5356 27829 5365 27863
rect 5365 27829 5399 27863
rect 5399 27829 5408 27863
rect 5356 27820 5408 27829
rect 6092 27820 6144 27872
rect 7840 27863 7892 27872
rect 7840 27829 7849 27863
rect 7849 27829 7883 27863
rect 7883 27829 7892 27863
rect 7840 27820 7892 27829
rect 19340 27888 19392 27940
rect 21824 27888 21876 27940
rect 11152 27863 11204 27872
rect 11152 27829 11161 27863
rect 11161 27829 11195 27863
rect 11195 27829 11204 27863
rect 11152 27820 11204 27829
rect 11612 27820 11664 27872
rect 20720 27820 20772 27872
rect 23480 27888 23532 27940
rect 23020 27820 23072 27872
rect 23756 27999 23808 28008
rect 23756 27965 23765 27999
rect 23765 27965 23799 27999
rect 23799 27965 23808 27999
rect 23756 27956 23808 27965
rect 24032 27863 24084 27872
rect 24032 27829 24041 27863
rect 24041 27829 24075 27863
rect 24075 27829 24084 27863
rect 24032 27820 24084 27829
rect 4182 27718 4234 27770
rect 4246 27718 4298 27770
rect 4310 27718 4362 27770
rect 4374 27718 4426 27770
rect 4438 27718 4490 27770
rect 4502 27718 4554 27770
rect 10182 27718 10234 27770
rect 10246 27718 10298 27770
rect 10310 27718 10362 27770
rect 10374 27718 10426 27770
rect 10438 27718 10490 27770
rect 10502 27718 10554 27770
rect 16182 27718 16234 27770
rect 16246 27718 16298 27770
rect 16310 27718 16362 27770
rect 16374 27718 16426 27770
rect 16438 27718 16490 27770
rect 16502 27718 16554 27770
rect 22182 27718 22234 27770
rect 22246 27718 22298 27770
rect 22310 27718 22362 27770
rect 22374 27718 22426 27770
rect 22438 27718 22490 27770
rect 22502 27718 22554 27770
rect 28182 27718 28234 27770
rect 28246 27718 28298 27770
rect 28310 27718 28362 27770
rect 28374 27718 28426 27770
rect 28438 27718 28490 27770
rect 28502 27718 28554 27770
rect 4620 27616 4672 27668
rect 6460 27616 6512 27668
rect 7196 27616 7248 27668
rect 8760 27616 8812 27668
rect 9128 27616 9180 27668
rect 13636 27659 13688 27668
rect 13636 27625 13645 27659
rect 13645 27625 13679 27659
rect 13679 27625 13688 27659
rect 13636 27616 13688 27625
rect 15752 27616 15804 27668
rect 22008 27659 22060 27668
rect 22008 27625 22017 27659
rect 22017 27625 22051 27659
rect 22051 27625 22060 27659
rect 22008 27616 22060 27625
rect 22928 27616 22980 27668
rect 5356 27412 5408 27464
rect 7472 27548 7524 27600
rect 7840 27480 7892 27532
rect 13728 27548 13780 27600
rect 16580 27548 16632 27600
rect 22376 27548 22428 27600
rect 6092 27344 6144 27396
rect 7196 27455 7248 27464
rect 7196 27421 7205 27455
rect 7205 27421 7239 27455
rect 7239 27421 7248 27455
rect 7196 27412 7248 27421
rect 7656 27412 7708 27464
rect 7748 27412 7800 27464
rect 11980 27455 12032 27464
rect 11980 27421 11989 27455
rect 11989 27421 12023 27455
rect 12023 27421 12032 27455
rect 11980 27412 12032 27421
rect 12348 27412 12400 27464
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 6552 27319 6604 27328
rect 6552 27285 6561 27319
rect 6561 27285 6595 27319
rect 6595 27285 6604 27319
rect 6552 27276 6604 27285
rect 14096 27319 14148 27328
rect 14096 27285 14105 27319
rect 14105 27285 14139 27319
rect 14139 27285 14148 27319
rect 14096 27276 14148 27285
rect 16028 27276 16080 27328
rect 16580 27455 16632 27464
rect 16580 27421 16589 27455
rect 16589 27421 16623 27455
rect 16623 27421 16632 27455
rect 16580 27412 16632 27421
rect 20996 27523 21048 27532
rect 20996 27489 21005 27523
rect 21005 27489 21039 27523
rect 21039 27489 21048 27523
rect 20996 27480 21048 27489
rect 16672 27344 16724 27396
rect 19432 27412 19484 27464
rect 22652 27480 22704 27532
rect 21548 27455 21600 27464
rect 21548 27421 21557 27455
rect 21557 27421 21591 27455
rect 21591 27421 21600 27455
rect 21548 27412 21600 27421
rect 21916 27412 21968 27464
rect 22928 27480 22980 27532
rect 24860 27523 24912 27532
rect 24860 27489 24869 27523
rect 24869 27489 24903 27523
rect 24903 27489 24912 27523
rect 24860 27480 24912 27489
rect 16856 27276 16908 27328
rect 19708 27276 19760 27328
rect 20444 27319 20496 27328
rect 20444 27285 20453 27319
rect 20453 27285 20487 27319
rect 20487 27285 20496 27319
rect 20444 27276 20496 27285
rect 23388 27412 23440 27464
rect 24952 27412 25004 27464
rect 26148 27455 26200 27464
rect 26148 27421 26157 27455
rect 26157 27421 26191 27455
rect 26191 27421 26200 27455
rect 26148 27412 26200 27421
rect 22468 27276 22520 27328
rect 22560 27276 22612 27328
rect 26332 27276 26384 27328
rect 26700 27387 26752 27396
rect 26700 27353 26709 27387
rect 26709 27353 26743 27387
rect 26743 27353 26752 27387
rect 26700 27344 26752 27353
rect 27344 27344 27396 27396
rect 27252 27276 27304 27328
rect 4922 27174 4974 27226
rect 4986 27174 5038 27226
rect 5050 27174 5102 27226
rect 5114 27174 5166 27226
rect 5178 27174 5230 27226
rect 5242 27174 5294 27226
rect 10922 27174 10974 27226
rect 10986 27174 11038 27226
rect 11050 27174 11102 27226
rect 11114 27174 11166 27226
rect 11178 27174 11230 27226
rect 11242 27174 11294 27226
rect 16922 27174 16974 27226
rect 16986 27174 17038 27226
rect 17050 27174 17102 27226
rect 17114 27174 17166 27226
rect 17178 27174 17230 27226
rect 17242 27174 17294 27226
rect 22922 27174 22974 27226
rect 22986 27174 23038 27226
rect 23050 27174 23102 27226
rect 23114 27174 23166 27226
rect 23178 27174 23230 27226
rect 23242 27174 23294 27226
rect 28922 27174 28974 27226
rect 28986 27174 29038 27226
rect 29050 27174 29102 27226
rect 29114 27174 29166 27226
rect 29178 27174 29230 27226
rect 29242 27174 29294 27226
rect 11980 27072 12032 27124
rect 14096 27072 14148 27124
rect 15752 27072 15804 27124
rect 13176 27047 13228 27056
rect 13176 27013 13185 27047
rect 13185 27013 13219 27047
rect 13219 27013 13228 27047
rect 13176 27004 13228 27013
rect 16764 27004 16816 27056
rect 20444 27072 20496 27124
rect 21548 27072 21600 27124
rect 22008 27072 22060 27124
rect 22376 27072 22428 27124
rect 22468 27004 22520 27056
rect 17040 26868 17092 26920
rect 17316 26868 17368 26920
rect 19984 26868 20036 26920
rect 21824 26868 21876 26920
rect 22560 26868 22612 26920
rect 22652 26800 22704 26852
rect 10048 26775 10100 26784
rect 10048 26741 10057 26775
rect 10057 26741 10091 26775
rect 10091 26741 10100 26775
rect 10048 26732 10100 26741
rect 10692 26732 10744 26784
rect 13636 26732 13688 26784
rect 21364 26732 21416 26784
rect 23480 27072 23532 27124
rect 23756 27072 23808 27124
rect 26148 27072 26200 27124
rect 25780 27004 25832 27056
rect 26332 27072 26384 27124
rect 24400 26936 24452 26988
rect 24216 26868 24268 26920
rect 25044 26868 25096 26920
rect 24400 26800 24452 26852
rect 24768 26800 24820 26852
rect 23848 26732 23900 26784
rect 24492 26732 24544 26784
rect 4182 26630 4234 26682
rect 4246 26630 4298 26682
rect 4310 26630 4362 26682
rect 4374 26630 4426 26682
rect 4438 26630 4490 26682
rect 4502 26630 4554 26682
rect 10182 26630 10234 26682
rect 10246 26630 10298 26682
rect 10310 26630 10362 26682
rect 10374 26630 10426 26682
rect 10438 26630 10490 26682
rect 10502 26630 10554 26682
rect 16182 26630 16234 26682
rect 16246 26630 16298 26682
rect 16310 26630 16362 26682
rect 16374 26630 16426 26682
rect 16438 26630 16490 26682
rect 16502 26630 16554 26682
rect 22182 26630 22234 26682
rect 22246 26630 22298 26682
rect 22310 26630 22362 26682
rect 22374 26630 22426 26682
rect 22438 26630 22490 26682
rect 22502 26630 22554 26682
rect 28182 26630 28234 26682
rect 28246 26630 28298 26682
rect 28310 26630 28362 26682
rect 28374 26630 28426 26682
rect 28438 26630 28490 26682
rect 28502 26630 28554 26682
rect 11428 26528 11480 26580
rect 10692 26460 10744 26512
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 9588 26324 9640 26376
rect 10508 26324 10560 26376
rect 16672 26528 16724 26580
rect 19708 26528 19760 26580
rect 21824 26571 21876 26580
rect 21824 26537 21833 26571
rect 21833 26537 21867 26571
rect 21867 26537 21876 26571
rect 21824 26528 21876 26537
rect 13636 26460 13688 26512
rect 15200 26460 15252 26512
rect 15292 26392 15344 26444
rect 20260 26460 20312 26512
rect 16028 26392 16080 26444
rect 17040 26435 17092 26444
rect 17040 26401 17049 26435
rect 17049 26401 17083 26435
rect 17083 26401 17092 26435
rect 17040 26392 17092 26401
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 12440 26324 12492 26376
rect 14648 26367 14700 26376
rect 14648 26333 14657 26367
rect 14657 26333 14691 26367
rect 14691 26333 14700 26367
rect 14648 26324 14700 26333
rect 11796 26256 11848 26308
rect 12164 26256 12216 26308
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 19984 26324 20036 26376
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 25044 26528 25096 26580
rect 25780 26503 25832 26512
rect 25780 26469 25789 26503
rect 25789 26469 25823 26503
rect 25823 26469 25832 26503
rect 25780 26460 25832 26469
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 10416 26231 10468 26240
rect 10416 26197 10425 26231
rect 10425 26197 10459 26231
rect 10459 26197 10468 26231
rect 10416 26188 10468 26197
rect 11704 26231 11756 26240
rect 11704 26197 11713 26231
rect 11713 26197 11747 26231
rect 11747 26197 11756 26231
rect 11704 26188 11756 26197
rect 12900 26188 12952 26240
rect 21364 26256 21416 26308
rect 17960 26188 18012 26240
rect 4922 26086 4974 26138
rect 4986 26086 5038 26138
rect 5050 26086 5102 26138
rect 5114 26086 5166 26138
rect 5178 26086 5230 26138
rect 5242 26086 5294 26138
rect 10922 26086 10974 26138
rect 10986 26086 11038 26138
rect 11050 26086 11102 26138
rect 11114 26086 11166 26138
rect 11178 26086 11230 26138
rect 11242 26086 11294 26138
rect 16922 26086 16974 26138
rect 16986 26086 17038 26138
rect 17050 26086 17102 26138
rect 17114 26086 17166 26138
rect 17178 26086 17230 26138
rect 17242 26086 17294 26138
rect 22922 26086 22974 26138
rect 22986 26086 23038 26138
rect 23050 26086 23102 26138
rect 23114 26086 23166 26138
rect 23178 26086 23230 26138
rect 23242 26086 23294 26138
rect 28922 26086 28974 26138
rect 28986 26086 29038 26138
rect 29050 26086 29102 26138
rect 29114 26086 29166 26138
rect 29178 26086 29230 26138
rect 29242 26086 29294 26138
rect 8576 25984 8628 26036
rect 10048 25984 10100 26036
rect 10416 25984 10468 26036
rect 12900 25916 12952 25968
rect 14648 25984 14700 26036
rect 24032 25984 24084 26036
rect 19984 25959 20036 25968
rect 19984 25925 19993 25959
rect 19993 25925 20027 25959
rect 20027 25925 20036 25959
rect 19984 25916 20036 25925
rect 7380 25848 7432 25900
rect 8116 25891 8168 25900
rect 8116 25857 8150 25891
rect 8150 25857 8168 25891
rect 8116 25848 8168 25857
rect 9680 25848 9732 25900
rect 5540 25823 5592 25832
rect 5540 25789 5549 25823
rect 5549 25789 5583 25823
rect 5583 25789 5592 25823
rect 5540 25780 5592 25789
rect 12440 25848 12492 25900
rect 17960 25848 18012 25900
rect 25780 25848 25832 25900
rect 9956 25823 10008 25832
rect 9956 25789 9965 25823
rect 9965 25789 9999 25823
rect 9999 25789 10008 25823
rect 9956 25780 10008 25789
rect 10600 25780 10652 25832
rect 12348 25780 12400 25832
rect 12532 25780 12584 25832
rect 20260 25780 20312 25832
rect 24492 25780 24544 25832
rect 10508 25712 10560 25764
rect 24860 25780 24912 25832
rect 4896 25687 4948 25696
rect 4896 25653 4905 25687
rect 4905 25653 4939 25687
rect 4939 25653 4948 25687
rect 4896 25644 4948 25653
rect 7012 25644 7064 25696
rect 8852 25644 8904 25696
rect 9312 25644 9364 25696
rect 11980 25644 12032 25696
rect 13084 25644 13136 25696
rect 14740 25644 14792 25696
rect 4182 25542 4234 25594
rect 4246 25542 4298 25594
rect 4310 25542 4362 25594
rect 4374 25542 4426 25594
rect 4438 25542 4490 25594
rect 4502 25542 4554 25594
rect 10182 25542 10234 25594
rect 10246 25542 10298 25594
rect 10310 25542 10362 25594
rect 10374 25542 10426 25594
rect 10438 25542 10490 25594
rect 10502 25542 10554 25594
rect 16182 25542 16234 25594
rect 16246 25542 16298 25594
rect 16310 25542 16362 25594
rect 16374 25542 16426 25594
rect 16438 25542 16490 25594
rect 16502 25542 16554 25594
rect 22182 25542 22234 25594
rect 22246 25542 22298 25594
rect 22310 25542 22362 25594
rect 22374 25542 22426 25594
rect 22438 25542 22490 25594
rect 22502 25542 22554 25594
rect 28182 25542 28234 25594
rect 28246 25542 28298 25594
rect 28310 25542 28362 25594
rect 28374 25542 28426 25594
rect 28438 25542 28490 25594
rect 28502 25542 28554 25594
rect 4896 25440 4948 25492
rect 5356 25440 5408 25492
rect 6000 25440 6052 25492
rect 3976 25143 4028 25152
rect 3976 25109 3985 25143
rect 3985 25109 4019 25143
rect 4019 25109 4028 25143
rect 3976 25100 4028 25109
rect 4712 25236 4764 25288
rect 7380 25440 7432 25492
rect 8116 25440 8168 25492
rect 9312 25440 9364 25492
rect 9588 25440 9640 25492
rect 12348 25440 12400 25492
rect 6644 25372 6696 25424
rect 5448 25168 5500 25220
rect 6828 25168 6880 25220
rect 7472 25304 7524 25356
rect 31300 25372 31352 25424
rect 11612 25347 11664 25356
rect 11612 25313 11621 25347
rect 11621 25313 11655 25347
rect 11655 25313 11664 25347
rect 11612 25304 11664 25313
rect 17868 25304 17920 25356
rect 18880 25347 18932 25356
rect 18880 25313 18889 25347
rect 18889 25313 18923 25347
rect 18923 25313 18932 25347
rect 18880 25304 18932 25313
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 4804 25100 4856 25152
rect 6092 25100 6144 25152
rect 6920 25143 6972 25152
rect 6920 25109 6929 25143
rect 6929 25109 6963 25143
rect 6963 25109 6972 25143
rect 6920 25100 6972 25109
rect 12348 25211 12400 25220
rect 12348 25177 12382 25211
rect 12382 25177 12400 25211
rect 12348 25168 12400 25177
rect 18420 25168 18472 25220
rect 19800 25279 19852 25288
rect 19800 25245 19809 25279
rect 19809 25245 19843 25279
rect 19843 25245 19852 25279
rect 19800 25236 19852 25245
rect 30656 25279 30708 25288
rect 30656 25245 30665 25279
rect 30665 25245 30699 25279
rect 30699 25245 30708 25279
rect 30656 25236 30708 25245
rect 20812 25168 20864 25220
rect 9956 25100 10008 25152
rect 12532 25100 12584 25152
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 17500 25100 17552 25109
rect 18328 25143 18380 25152
rect 18328 25109 18337 25143
rect 18337 25109 18371 25143
rect 18371 25109 18380 25143
rect 18328 25100 18380 25109
rect 20628 25100 20680 25152
rect 4922 24998 4974 25050
rect 4986 24998 5038 25050
rect 5050 24998 5102 25050
rect 5114 24998 5166 25050
rect 5178 24998 5230 25050
rect 5242 24998 5294 25050
rect 10922 24998 10974 25050
rect 10986 24998 11038 25050
rect 11050 24998 11102 25050
rect 11114 24998 11166 25050
rect 11178 24998 11230 25050
rect 11242 24998 11294 25050
rect 16922 24998 16974 25050
rect 16986 24998 17038 25050
rect 17050 24998 17102 25050
rect 17114 24998 17166 25050
rect 17178 24998 17230 25050
rect 17242 24998 17294 25050
rect 22922 24998 22974 25050
rect 22986 24998 23038 25050
rect 23050 24998 23102 25050
rect 23114 24998 23166 25050
rect 23178 24998 23230 25050
rect 23242 24998 23294 25050
rect 28922 24998 28974 25050
rect 28986 24998 29038 25050
rect 29050 24998 29102 25050
rect 29114 24998 29166 25050
rect 29178 24998 29230 25050
rect 29242 24998 29294 25050
rect 4712 24896 4764 24948
rect 5448 24939 5500 24948
rect 5448 24905 5457 24939
rect 5457 24905 5491 24939
rect 5491 24905 5500 24939
rect 5448 24896 5500 24905
rect 4804 24828 4856 24880
rect 3976 24803 4028 24812
rect 3976 24769 4010 24803
rect 4010 24769 4028 24803
rect 6092 24828 6144 24880
rect 6644 24871 6696 24880
rect 6644 24837 6653 24871
rect 6653 24837 6687 24871
rect 6687 24837 6696 24871
rect 6644 24828 6696 24837
rect 7380 24828 7432 24880
rect 8116 24871 8168 24880
rect 8116 24837 8125 24871
rect 8125 24837 8159 24871
rect 8159 24837 8168 24871
rect 8116 24828 8168 24837
rect 9312 24896 9364 24948
rect 9956 24939 10008 24948
rect 9956 24905 9965 24939
rect 9965 24905 9999 24939
rect 9999 24905 10008 24939
rect 9956 24896 10008 24905
rect 12348 24896 12400 24948
rect 12440 24896 12492 24948
rect 9680 24828 9732 24880
rect 12532 24828 12584 24880
rect 3976 24760 4028 24769
rect 5540 24624 5592 24676
rect 7656 24760 7708 24812
rect 10692 24760 10744 24812
rect 11612 24760 11664 24812
rect 7196 24692 7248 24744
rect 9680 24692 9732 24744
rect 10140 24735 10192 24744
rect 10140 24701 10149 24735
rect 10149 24701 10183 24735
rect 10183 24701 10192 24735
rect 10140 24692 10192 24701
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 11428 24556 11480 24608
rect 12164 24760 12216 24812
rect 14096 24896 14148 24948
rect 14648 24896 14700 24948
rect 17500 24896 17552 24948
rect 18420 24896 18472 24948
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 19616 24828 19668 24880
rect 17592 24760 17644 24812
rect 11980 24556 12032 24608
rect 12072 24599 12124 24608
rect 12072 24565 12081 24599
rect 12081 24565 12115 24599
rect 12115 24565 12124 24599
rect 12072 24556 12124 24565
rect 13452 24624 13504 24676
rect 13360 24599 13412 24608
rect 13360 24565 13369 24599
rect 13369 24565 13403 24599
rect 13403 24565 13412 24599
rect 13360 24556 13412 24565
rect 14556 24692 14608 24744
rect 14924 24735 14976 24744
rect 14924 24701 14933 24735
rect 14933 24701 14967 24735
rect 14967 24701 14976 24735
rect 14924 24692 14976 24701
rect 13728 24624 13780 24676
rect 19800 24692 19852 24744
rect 20352 24760 20404 24812
rect 20812 24803 20864 24812
rect 20812 24769 20821 24803
rect 20821 24769 20855 24803
rect 20855 24769 20864 24803
rect 20812 24760 20864 24769
rect 21364 24803 21416 24812
rect 21364 24769 21373 24803
rect 21373 24769 21407 24803
rect 21407 24769 21416 24803
rect 21364 24760 21416 24769
rect 14372 24599 14424 24608
rect 14372 24565 14381 24599
rect 14381 24565 14415 24599
rect 14415 24565 14424 24599
rect 14372 24556 14424 24565
rect 17224 24599 17276 24608
rect 17224 24565 17233 24599
rect 17233 24565 17267 24599
rect 17267 24565 17276 24599
rect 17224 24556 17276 24565
rect 17500 24556 17552 24608
rect 18420 24556 18472 24608
rect 19892 24624 19944 24676
rect 20904 24735 20956 24744
rect 20904 24701 20913 24735
rect 20913 24701 20947 24735
rect 20947 24701 20956 24735
rect 20904 24692 20956 24701
rect 21272 24692 21324 24744
rect 24400 24735 24452 24744
rect 24400 24701 24409 24735
rect 24409 24701 24443 24735
rect 24443 24701 24452 24735
rect 24400 24692 24452 24701
rect 25228 24735 25280 24744
rect 25228 24701 25237 24735
rect 25237 24701 25271 24735
rect 25271 24701 25280 24735
rect 25228 24692 25280 24701
rect 23572 24624 23624 24676
rect 20260 24599 20312 24608
rect 20260 24565 20269 24599
rect 20269 24565 20303 24599
rect 20303 24565 20312 24599
rect 20260 24556 20312 24565
rect 21180 24599 21232 24608
rect 21180 24565 21189 24599
rect 21189 24565 21223 24599
rect 21223 24565 21232 24599
rect 21180 24556 21232 24565
rect 22100 24556 22152 24608
rect 24676 24624 24728 24676
rect 23848 24599 23900 24608
rect 23848 24565 23857 24599
rect 23857 24565 23891 24599
rect 23891 24565 23900 24599
rect 23848 24556 23900 24565
rect 24584 24599 24636 24608
rect 24584 24565 24593 24599
rect 24593 24565 24627 24599
rect 24627 24565 24636 24599
rect 24584 24556 24636 24565
rect 4182 24454 4234 24506
rect 4246 24454 4298 24506
rect 4310 24454 4362 24506
rect 4374 24454 4426 24506
rect 4438 24454 4490 24506
rect 4502 24454 4554 24506
rect 10182 24454 10234 24506
rect 10246 24454 10298 24506
rect 10310 24454 10362 24506
rect 10374 24454 10426 24506
rect 10438 24454 10490 24506
rect 10502 24454 10554 24506
rect 16182 24454 16234 24506
rect 16246 24454 16298 24506
rect 16310 24454 16362 24506
rect 16374 24454 16426 24506
rect 16438 24454 16490 24506
rect 16502 24454 16554 24506
rect 22182 24454 22234 24506
rect 22246 24454 22298 24506
rect 22310 24454 22362 24506
rect 22374 24454 22426 24506
rect 22438 24454 22490 24506
rect 22502 24454 22554 24506
rect 28182 24454 28234 24506
rect 28246 24454 28298 24506
rect 28310 24454 28362 24506
rect 28374 24454 28426 24506
rect 28438 24454 28490 24506
rect 28502 24454 28554 24506
rect 6920 24352 6972 24404
rect 12072 24352 12124 24404
rect 8576 24191 8628 24200
rect 8576 24157 8585 24191
rect 8585 24157 8619 24191
rect 8619 24157 8628 24191
rect 8576 24148 8628 24157
rect 10784 24148 10836 24200
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 13360 24352 13412 24404
rect 14924 24352 14976 24404
rect 18420 24395 18472 24404
rect 18420 24361 18429 24395
rect 18429 24361 18463 24395
rect 18463 24361 18472 24395
rect 18420 24352 18472 24361
rect 19892 24352 19944 24404
rect 20168 24352 20220 24404
rect 16120 24216 16172 24268
rect 21272 24395 21324 24404
rect 21272 24361 21281 24395
rect 21281 24361 21315 24395
rect 21315 24361 21324 24395
rect 21272 24352 21324 24361
rect 21364 24395 21416 24404
rect 21364 24361 21373 24395
rect 21373 24361 21407 24395
rect 21407 24361 21416 24395
rect 21364 24352 21416 24361
rect 22100 24284 22152 24336
rect 15108 24148 15160 24200
rect 20996 24216 21048 24268
rect 940 24080 992 24132
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 13820 24080 13872 24132
rect 8392 24055 8444 24064
rect 8392 24021 8401 24055
rect 8401 24021 8435 24055
rect 8435 24021 8444 24055
rect 8392 24012 8444 24021
rect 9680 24055 9732 24064
rect 9680 24021 9689 24055
rect 9689 24021 9723 24055
rect 9723 24021 9732 24055
rect 9680 24012 9732 24021
rect 12256 24012 12308 24064
rect 13728 24012 13780 24064
rect 15292 24012 15344 24064
rect 15752 24055 15804 24064
rect 15752 24021 15761 24055
rect 15761 24021 15795 24055
rect 15795 24021 15804 24055
rect 15752 24012 15804 24021
rect 17224 24080 17276 24132
rect 17500 24080 17552 24132
rect 20444 24148 20496 24200
rect 20628 24148 20680 24200
rect 24400 24352 24452 24404
rect 24584 24352 24636 24404
rect 24860 24352 24912 24404
rect 19984 24080 20036 24132
rect 23756 24148 23808 24200
rect 24676 24216 24728 24268
rect 21824 24055 21876 24064
rect 21824 24021 21833 24055
rect 21833 24021 21867 24055
rect 21867 24021 21876 24055
rect 21824 24012 21876 24021
rect 22836 24012 22888 24064
rect 24124 24012 24176 24064
rect 25596 24055 25648 24064
rect 25596 24021 25605 24055
rect 25605 24021 25639 24055
rect 25639 24021 25648 24055
rect 25596 24012 25648 24021
rect 25964 24055 26016 24064
rect 25964 24021 25973 24055
rect 25973 24021 26007 24055
rect 26007 24021 26016 24055
rect 25964 24012 26016 24021
rect 26884 24012 26936 24064
rect 4922 23910 4974 23962
rect 4986 23910 5038 23962
rect 5050 23910 5102 23962
rect 5114 23910 5166 23962
rect 5178 23910 5230 23962
rect 5242 23910 5294 23962
rect 10922 23910 10974 23962
rect 10986 23910 11038 23962
rect 11050 23910 11102 23962
rect 11114 23910 11166 23962
rect 11178 23910 11230 23962
rect 11242 23910 11294 23962
rect 16922 23910 16974 23962
rect 16986 23910 17038 23962
rect 17050 23910 17102 23962
rect 17114 23910 17166 23962
rect 17178 23910 17230 23962
rect 17242 23910 17294 23962
rect 22922 23910 22974 23962
rect 22986 23910 23038 23962
rect 23050 23910 23102 23962
rect 23114 23910 23166 23962
rect 23178 23910 23230 23962
rect 23242 23910 23294 23962
rect 28922 23910 28974 23962
rect 28986 23910 29038 23962
rect 29050 23910 29102 23962
rect 29114 23910 29166 23962
rect 29178 23910 29230 23962
rect 29242 23910 29294 23962
rect 8392 23808 8444 23860
rect 8576 23808 8628 23860
rect 9680 23808 9732 23860
rect 13452 23808 13504 23860
rect 13728 23808 13780 23860
rect 13820 23851 13872 23860
rect 13820 23817 13829 23851
rect 13829 23817 13863 23851
rect 13863 23817 13872 23851
rect 13820 23808 13872 23817
rect 8116 23672 8168 23724
rect 9956 23715 10008 23724
rect 9956 23681 9965 23715
rect 9965 23681 9999 23715
rect 9999 23681 10008 23715
rect 9956 23672 10008 23681
rect 4620 23511 4672 23520
rect 4620 23477 4629 23511
rect 4629 23477 4663 23511
rect 4663 23477 4672 23511
rect 4620 23468 4672 23477
rect 5356 23604 5408 23656
rect 5908 23604 5960 23656
rect 6000 23647 6052 23656
rect 6000 23613 6009 23647
rect 6009 23613 6043 23647
rect 6043 23613 6052 23647
rect 6000 23604 6052 23613
rect 9864 23604 9916 23656
rect 10784 23536 10836 23588
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 13452 23672 13504 23724
rect 13544 23672 13596 23724
rect 14372 23808 14424 23860
rect 15108 23808 15160 23860
rect 16120 23808 16172 23860
rect 17592 23851 17644 23860
rect 17592 23817 17601 23851
rect 17601 23817 17635 23851
rect 17635 23817 17644 23851
rect 17592 23808 17644 23817
rect 18328 23808 18380 23860
rect 20260 23808 20312 23860
rect 21180 23808 21232 23860
rect 21824 23851 21876 23860
rect 21824 23817 21833 23851
rect 21833 23817 21867 23851
rect 21867 23817 21876 23851
rect 21824 23808 21876 23817
rect 23848 23808 23900 23860
rect 24124 23808 24176 23860
rect 17868 23783 17920 23792
rect 17868 23749 17877 23783
rect 17877 23749 17911 23783
rect 17911 23749 17920 23783
rect 17868 23740 17920 23749
rect 13912 23604 13964 23656
rect 13452 23536 13504 23588
rect 14556 23647 14608 23656
rect 14556 23613 14565 23647
rect 14565 23613 14599 23647
rect 14599 23613 14608 23647
rect 14556 23604 14608 23613
rect 16212 23672 16264 23724
rect 17224 23672 17276 23724
rect 19984 23672 20036 23724
rect 22652 23740 22704 23792
rect 23756 23740 23808 23792
rect 9220 23468 9272 23520
rect 9772 23468 9824 23520
rect 10600 23468 10652 23520
rect 12440 23468 12492 23520
rect 18880 23468 18932 23520
rect 20260 23468 20312 23520
rect 20996 23468 21048 23520
rect 23480 23672 23532 23724
rect 23572 23715 23624 23724
rect 23572 23681 23581 23715
rect 23581 23681 23615 23715
rect 23615 23681 23624 23715
rect 23572 23672 23624 23681
rect 22100 23536 22152 23588
rect 23664 23647 23716 23656
rect 23664 23613 23673 23647
rect 23673 23613 23707 23647
rect 23707 23613 23716 23647
rect 23664 23604 23716 23613
rect 23848 23604 23900 23656
rect 25596 23808 25648 23860
rect 25964 23808 26016 23860
rect 24124 23604 24176 23656
rect 26332 23647 26384 23656
rect 26332 23613 26341 23647
rect 26341 23613 26375 23647
rect 26375 23613 26384 23647
rect 26332 23604 26384 23613
rect 23020 23511 23072 23520
rect 23020 23477 23029 23511
rect 23029 23477 23063 23511
rect 23063 23477 23072 23511
rect 23020 23468 23072 23477
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 23756 23468 23808 23520
rect 25228 23468 25280 23520
rect 26516 23511 26568 23520
rect 26516 23477 26525 23511
rect 26525 23477 26559 23511
rect 26559 23477 26568 23511
rect 26516 23468 26568 23477
rect 4182 23366 4234 23418
rect 4246 23366 4298 23418
rect 4310 23366 4362 23418
rect 4374 23366 4426 23418
rect 4438 23366 4490 23418
rect 4502 23366 4554 23418
rect 10182 23366 10234 23418
rect 10246 23366 10298 23418
rect 10310 23366 10362 23418
rect 10374 23366 10426 23418
rect 10438 23366 10490 23418
rect 10502 23366 10554 23418
rect 16182 23366 16234 23418
rect 16246 23366 16298 23418
rect 16310 23366 16362 23418
rect 16374 23366 16426 23418
rect 16438 23366 16490 23418
rect 16502 23366 16554 23418
rect 22182 23366 22234 23418
rect 22246 23366 22298 23418
rect 22310 23366 22362 23418
rect 22374 23366 22426 23418
rect 22438 23366 22490 23418
rect 22502 23366 22554 23418
rect 28182 23366 28234 23418
rect 28246 23366 28298 23418
rect 28310 23366 28362 23418
rect 28374 23366 28426 23418
rect 28438 23366 28490 23418
rect 28502 23366 28554 23418
rect 4712 23264 4764 23316
rect 4620 23060 4672 23112
rect 7012 23264 7064 23316
rect 9956 23264 10008 23316
rect 10876 23264 10928 23316
rect 11520 23264 11572 23316
rect 13912 23307 13964 23316
rect 13912 23273 13921 23307
rect 13921 23273 13955 23307
rect 13955 23273 13964 23307
rect 13912 23264 13964 23273
rect 16028 23264 16080 23316
rect 22652 23264 22704 23316
rect 22836 23264 22888 23316
rect 23480 23264 23532 23316
rect 24492 23307 24544 23316
rect 24492 23273 24501 23307
rect 24501 23273 24535 23307
rect 24535 23273 24544 23307
rect 24492 23264 24544 23273
rect 26332 23264 26384 23316
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 9220 23128 9272 23180
rect 8116 23060 8168 23112
rect 9772 23128 9824 23180
rect 11888 23196 11940 23248
rect 9864 23060 9916 23112
rect 10232 23060 10284 23112
rect 10600 23060 10652 23112
rect 11704 23128 11756 23180
rect 12440 23128 12492 23180
rect 12532 23171 12584 23180
rect 12532 23137 12541 23171
rect 12541 23137 12575 23171
rect 12575 23137 12584 23171
rect 12532 23128 12584 23137
rect 15476 23128 15528 23180
rect 17776 23128 17828 23180
rect 20444 23128 20496 23180
rect 24124 23128 24176 23180
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 10876 23060 10928 23069
rect 12256 23103 12308 23112
rect 12256 23069 12265 23103
rect 12265 23069 12299 23103
rect 12299 23069 12308 23103
rect 12256 23060 12308 23069
rect 12624 23060 12676 23112
rect 15752 23060 15804 23112
rect 19340 23060 19392 23112
rect 21272 23060 21324 23112
rect 22100 23103 22152 23112
rect 22100 23069 22109 23103
rect 22109 23069 22143 23103
rect 22143 23069 22152 23103
rect 22100 23060 22152 23069
rect 22652 23060 22704 23112
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 5356 22992 5408 23044
rect 7748 22992 7800 23044
rect 11612 23035 11664 23044
rect 11612 23001 11621 23035
rect 11621 23001 11655 23035
rect 11655 23001 11664 23035
rect 11612 22992 11664 23001
rect 4252 22967 4304 22976
rect 4252 22933 4261 22967
rect 4261 22933 4295 22967
rect 4295 22933 4304 22967
rect 4252 22924 4304 22933
rect 6184 22967 6236 22976
rect 6184 22933 6193 22967
rect 6193 22933 6227 22967
rect 6227 22933 6236 22967
rect 6184 22924 6236 22933
rect 6276 22967 6328 22976
rect 6276 22933 6285 22967
rect 6285 22933 6319 22967
rect 6319 22933 6328 22967
rect 6276 22924 6328 22933
rect 6736 22967 6788 22976
rect 6736 22933 6745 22967
rect 6745 22933 6779 22967
rect 6779 22933 6788 22967
rect 6736 22924 6788 22933
rect 8944 22967 8996 22976
rect 8944 22933 8953 22967
rect 8953 22933 8987 22967
rect 8987 22933 8996 22967
rect 8944 22924 8996 22933
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 23296 22992 23348 23044
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 21824 22924 21876 22976
rect 24032 23035 24084 23044
rect 24032 23001 24041 23035
rect 24041 23001 24075 23035
rect 24075 23001 24084 23035
rect 24032 22992 24084 23001
rect 24400 23060 24452 23112
rect 25044 23060 25096 23112
rect 26516 23060 26568 23112
rect 25228 22992 25280 23044
rect 24400 22924 24452 22976
rect 4922 22822 4974 22874
rect 4986 22822 5038 22874
rect 5050 22822 5102 22874
rect 5114 22822 5166 22874
rect 5178 22822 5230 22874
rect 5242 22822 5294 22874
rect 10922 22822 10974 22874
rect 10986 22822 11038 22874
rect 11050 22822 11102 22874
rect 11114 22822 11166 22874
rect 11178 22822 11230 22874
rect 11242 22822 11294 22874
rect 16922 22822 16974 22874
rect 16986 22822 17038 22874
rect 17050 22822 17102 22874
rect 17114 22822 17166 22874
rect 17178 22822 17230 22874
rect 17242 22822 17294 22874
rect 22922 22822 22974 22874
rect 22986 22822 23038 22874
rect 23050 22822 23102 22874
rect 23114 22822 23166 22874
rect 23178 22822 23230 22874
rect 23242 22822 23294 22874
rect 28922 22822 28974 22874
rect 28986 22822 29038 22874
rect 29050 22822 29102 22874
rect 29114 22822 29166 22874
rect 29178 22822 29230 22874
rect 29242 22822 29294 22874
rect 4252 22720 4304 22772
rect 5356 22763 5408 22772
rect 5356 22729 5365 22763
rect 5365 22729 5399 22763
rect 5399 22729 5408 22763
rect 5356 22720 5408 22729
rect 6276 22720 6328 22772
rect 6736 22720 6788 22772
rect 7196 22720 7248 22772
rect 7748 22720 7800 22772
rect 8944 22720 8996 22772
rect 11612 22720 11664 22772
rect 12256 22720 12308 22772
rect 14096 22720 14148 22772
rect 6368 22584 6420 22636
rect 3884 22559 3936 22568
rect 3884 22525 3893 22559
rect 3893 22525 3927 22559
rect 3927 22525 3936 22559
rect 3884 22516 3936 22525
rect 6184 22516 6236 22568
rect 7656 22584 7708 22636
rect 6000 22448 6052 22500
rect 6368 22448 6420 22500
rect 11888 22652 11940 22704
rect 14924 22720 14976 22772
rect 23756 22763 23808 22772
rect 23756 22729 23765 22763
rect 23765 22729 23799 22763
rect 23799 22729 23808 22763
rect 23756 22720 23808 22729
rect 24492 22720 24544 22772
rect 14740 22695 14792 22704
rect 14740 22661 14749 22695
rect 14749 22661 14783 22695
rect 14783 22661 14792 22695
rect 14740 22652 14792 22661
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 14464 22584 14516 22636
rect 15108 22584 15160 22636
rect 23940 22627 23992 22636
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 13728 22516 13780 22568
rect 15200 22516 15252 22568
rect 24124 22516 24176 22568
rect 24768 22584 24820 22636
rect 12900 22448 12952 22500
rect 16764 22448 16816 22500
rect 23664 22448 23716 22500
rect 16948 22380 17000 22432
rect 18328 22380 18380 22432
rect 4182 22278 4234 22330
rect 4246 22278 4298 22330
rect 4310 22278 4362 22330
rect 4374 22278 4426 22330
rect 4438 22278 4490 22330
rect 4502 22278 4554 22330
rect 10182 22278 10234 22330
rect 10246 22278 10298 22330
rect 10310 22278 10362 22330
rect 10374 22278 10426 22330
rect 10438 22278 10490 22330
rect 10502 22278 10554 22330
rect 16182 22278 16234 22330
rect 16246 22278 16298 22330
rect 16310 22278 16362 22330
rect 16374 22278 16426 22330
rect 16438 22278 16490 22330
rect 16502 22278 16554 22330
rect 22182 22278 22234 22330
rect 22246 22278 22298 22330
rect 22310 22278 22362 22330
rect 22374 22278 22426 22330
rect 22438 22278 22490 22330
rect 22502 22278 22554 22330
rect 28182 22278 28234 22330
rect 28246 22278 28298 22330
rect 28310 22278 28362 22330
rect 28374 22278 28426 22330
rect 28438 22278 28490 22330
rect 28502 22278 28554 22330
rect 9772 22176 9824 22228
rect 15200 22176 15252 22228
rect 15476 22176 15528 22228
rect 5724 22040 5776 22092
rect 8116 22040 8168 22092
rect 10784 22108 10836 22160
rect 11520 22108 11572 22160
rect 12900 22108 12952 22160
rect 14096 22151 14148 22160
rect 14096 22117 14105 22151
rect 14105 22117 14139 22151
rect 14139 22117 14148 22151
rect 14096 22108 14148 22117
rect 16580 22108 16632 22160
rect 7380 21972 7432 22024
rect 13268 22040 13320 22092
rect 17592 22108 17644 22160
rect 18880 22040 18932 22092
rect 9312 22015 9364 22024
rect 9312 21981 9321 22015
rect 9321 21981 9355 22015
rect 9355 21981 9364 22015
rect 9312 21972 9364 21981
rect 13084 21972 13136 22024
rect 11980 21904 12032 21956
rect 14464 21904 14516 21956
rect 7656 21836 7708 21888
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 8208 21836 8260 21845
rect 9680 21836 9732 21888
rect 9772 21836 9824 21888
rect 11612 21836 11664 21888
rect 11796 21836 11848 21888
rect 15844 21879 15896 21888
rect 15844 21845 15853 21879
rect 15853 21845 15887 21879
rect 15887 21845 15896 21879
rect 15844 21836 15896 21845
rect 16120 21904 16172 21956
rect 16304 21947 16356 21956
rect 16304 21913 16313 21947
rect 16313 21913 16347 21947
rect 16347 21913 16356 21947
rect 16304 21904 16356 21913
rect 16488 21947 16540 21956
rect 16488 21913 16497 21947
rect 16497 21913 16531 21947
rect 16531 21913 16540 21947
rect 16488 21904 16540 21913
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 24400 22151 24452 22160
rect 24400 22117 24409 22151
rect 24409 22117 24443 22151
rect 24443 22117 24452 22151
rect 24400 22108 24452 22117
rect 20536 22040 20588 22092
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 19432 21904 19484 21956
rect 19800 21904 19852 21956
rect 20168 21904 20220 21956
rect 20996 21879 21048 21888
rect 20996 21845 21005 21879
rect 21005 21845 21039 21879
rect 21039 21845 21048 21879
rect 20996 21836 21048 21845
rect 24032 21904 24084 21956
rect 24308 21904 24360 21956
rect 4922 21734 4974 21786
rect 4986 21734 5038 21786
rect 5050 21734 5102 21786
rect 5114 21734 5166 21786
rect 5178 21734 5230 21786
rect 5242 21734 5294 21786
rect 10922 21734 10974 21786
rect 10986 21734 11038 21786
rect 11050 21734 11102 21786
rect 11114 21734 11166 21786
rect 11178 21734 11230 21786
rect 11242 21734 11294 21786
rect 16922 21734 16974 21786
rect 16986 21734 17038 21786
rect 17050 21734 17102 21786
rect 17114 21734 17166 21786
rect 17178 21734 17230 21786
rect 17242 21734 17294 21786
rect 22922 21734 22974 21786
rect 22986 21734 23038 21786
rect 23050 21734 23102 21786
rect 23114 21734 23166 21786
rect 23178 21734 23230 21786
rect 23242 21734 23294 21786
rect 28922 21734 28974 21786
rect 28986 21734 29038 21786
rect 29050 21734 29102 21786
rect 29114 21734 29166 21786
rect 29178 21734 29230 21786
rect 29242 21734 29294 21786
rect 8208 21632 8260 21684
rect 10048 21632 10100 21684
rect 7380 21564 7432 21616
rect 13084 21675 13136 21684
rect 13084 21641 13093 21675
rect 13093 21641 13127 21675
rect 13127 21641 13136 21675
rect 13084 21632 13136 21641
rect 14096 21632 14148 21684
rect 15844 21632 15896 21684
rect 17408 21632 17460 21684
rect 20352 21632 20404 21684
rect 15200 21564 15252 21616
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 7564 21496 7616 21548
rect 9680 21496 9732 21548
rect 10692 21496 10744 21548
rect 12532 21496 12584 21548
rect 16948 21564 17000 21616
rect 18052 21564 18104 21616
rect 21824 21607 21876 21616
rect 21824 21573 21833 21607
rect 21833 21573 21867 21607
rect 21867 21573 21876 21607
rect 21824 21564 21876 21573
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 17132 21496 17184 21548
rect 7104 21428 7156 21480
rect 8760 21428 8812 21480
rect 5172 21292 5224 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 8300 21292 8352 21344
rect 8392 21292 8444 21344
rect 11060 21428 11112 21480
rect 11704 21471 11756 21480
rect 11704 21437 11713 21471
rect 11713 21437 11747 21471
rect 11747 21437 11756 21471
rect 11704 21428 11756 21437
rect 12992 21428 13044 21480
rect 13636 21471 13688 21480
rect 13636 21437 13645 21471
rect 13645 21437 13679 21471
rect 13679 21437 13688 21471
rect 13636 21428 13688 21437
rect 14556 21428 14608 21480
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 15844 21428 15896 21437
rect 16488 21471 16540 21480
rect 16488 21437 16497 21471
rect 16497 21437 16531 21471
rect 16531 21437 16540 21471
rect 16488 21428 16540 21437
rect 17224 21428 17276 21480
rect 9956 21292 10008 21344
rect 11612 21292 11664 21344
rect 13176 21335 13228 21344
rect 13176 21301 13185 21335
rect 13185 21301 13219 21335
rect 13219 21301 13228 21335
rect 13176 21292 13228 21301
rect 14740 21292 14792 21344
rect 16488 21292 16540 21344
rect 17868 21496 17920 21548
rect 22100 21496 22152 21548
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 17776 21471 17828 21480
rect 17776 21437 17785 21471
rect 17785 21437 17819 21471
rect 17819 21437 17828 21471
rect 17776 21428 17828 21437
rect 20904 21428 20956 21480
rect 23480 21428 23532 21480
rect 24032 21428 24084 21480
rect 24216 21539 24268 21548
rect 24216 21505 24225 21539
rect 24225 21505 24259 21539
rect 24259 21505 24268 21539
rect 24216 21496 24268 21505
rect 24216 21292 24268 21344
rect 24308 21335 24360 21344
rect 24308 21301 24317 21335
rect 24317 21301 24351 21335
rect 24351 21301 24360 21335
rect 24308 21292 24360 21301
rect 24400 21292 24452 21344
rect 4182 21190 4234 21242
rect 4246 21190 4298 21242
rect 4310 21190 4362 21242
rect 4374 21190 4426 21242
rect 4438 21190 4490 21242
rect 4502 21190 4554 21242
rect 10182 21190 10234 21242
rect 10246 21190 10298 21242
rect 10310 21190 10362 21242
rect 10374 21190 10426 21242
rect 10438 21190 10490 21242
rect 10502 21190 10554 21242
rect 16182 21190 16234 21242
rect 16246 21190 16298 21242
rect 16310 21190 16362 21242
rect 16374 21190 16426 21242
rect 16438 21190 16490 21242
rect 16502 21190 16554 21242
rect 22182 21190 22234 21242
rect 22246 21190 22298 21242
rect 22310 21190 22362 21242
rect 22374 21190 22426 21242
rect 22438 21190 22490 21242
rect 22502 21190 22554 21242
rect 28182 21190 28234 21242
rect 28246 21190 28298 21242
rect 28310 21190 28362 21242
rect 28374 21190 28426 21242
rect 28438 21190 28490 21242
rect 28502 21190 28554 21242
rect 5172 21131 5224 21140
rect 5172 21097 5181 21131
rect 5181 21097 5215 21131
rect 5215 21097 5224 21131
rect 5172 21088 5224 21097
rect 5448 21088 5500 21140
rect 3884 20884 3936 20936
rect 5908 20995 5960 21004
rect 5908 20961 5917 20995
rect 5917 20961 5951 20995
rect 5951 20961 5960 20995
rect 8392 21131 8444 21140
rect 8392 21097 8401 21131
rect 8401 21097 8435 21131
rect 8435 21097 8444 21131
rect 8392 21088 8444 21097
rect 9312 21088 9364 21140
rect 12532 21131 12584 21140
rect 12532 21097 12541 21131
rect 12541 21097 12575 21131
rect 12575 21097 12584 21131
rect 12532 21088 12584 21097
rect 13084 21088 13136 21140
rect 13176 21088 13228 21140
rect 13268 21088 13320 21140
rect 17224 21088 17276 21140
rect 17868 21088 17920 21140
rect 19340 21088 19392 21140
rect 19984 21088 20036 21140
rect 20168 21131 20220 21140
rect 20168 21097 20177 21131
rect 20177 21097 20211 21131
rect 20211 21097 20220 21131
rect 20168 21088 20220 21097
rect 22100 21088 22152 21140
rect 23756 21088 23808 21140
rect 23940 21088 23992 21140
rect 12992 21020 13044 21072
rect 5908 20952 5960 20961
rect 6644 20952 6696 21004
rect 8116 20952 8168 21004
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 4160 20816 4212 20868
rect 4804 20816 4856 20868
rect 7104 20884 7156 20936
rect 9680 20884 9732 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 10692 20884 10744 20936
rect 11428 20884 11480 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 12624 20884 12676 20936
rect 15844 21020 15896 21072
rect 13728 20952 13780 21004
rect 14648 20927 14700 20936
rect 14648 20893 14657 20927
rect 14657 20893 14691 20927
rect 14691 20893 14700 20927
rect 14648 20884 14700 20893
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 7472 20816 7524 20868
rect 11060 20816 11112 20868
rect 15292 20816 15344 20868
rect 16672 20952 16724 21004
rect 16764 20995 16816 21004
rect 16764 20961 16773 20995
rect 16773 20961 16807 20995
rect 16807 20961 16816 20995
rect 16764 20952 16816 20961
rect 16948 20952 17000 21004
rect 17500 20952 17552 21004
rect 24308 21020 24360 21072
rect 19616 20952 19668 21004
rect 16488 20884 16540 20936
rect 17684 20927 17736 20936
rect 17684 20893 17693 20927
rect 17693 20893 17727 20927
rect 17727 20893 17736 20927
rect 17684 20884 17736 20893
rect 18052 20884 18104 20936
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 20996 20884 21048 20936
rect 22468 20952 22520 21004
rect 23388 20952 23440 21004
rect 23480 20952 23532 21004
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 21732 20927 21784 20936
rect 21732 20893 21741 20927
rect 21741 20893 21775 20927
rect 21775 20893 21784 20927
rect 21732 20884 21784 20893
rect 18236 20816 18288 20868
rect 18328 20859 18380 20868
rect 18328 20825 18337 20859
rect 18337 20825 18371 20859
rect 18371 20825 18380 20859
rect 18328 20816 18380 20825
rect 5356 20748 5408 20800
rect 5724 20791 5776 20800
rect 5724 20757 5733 20791
rect 5733 20757 5767 20791
rect 5767 20757 5776 20791
rect 5724 20748 5776 20757
rect 6920 20791 6972 20800
rect 6920 20757 6929 20791
rect 6929 20757 6963 20791
rect 6963 20757 6972 20791
rect 6920 20748 6972 20757
rect 8484 20748 8536 20800
rect 8760 20748 8812 20800
rect 11428 20748 11480 20800
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 14096 20791 14148 20800
rect 14096 20757 14105 20791
rect 14105 20757 14139 20791
rect 14139 20757 14148 20791
rect 14096 20748 14148 20757
rect 17132 20748 17184 20800
rect 17684 20748 17736 20800
rect 19064 20816 19116 20868
rect 23756 20884 23808 20936
rect 23940 20927 23992 20936
rect 23940 20893 23949 20927
rect 23949 20893 23983 20927
rect 23983 20893 23992 20927
rect 23940 20884 23992 20893
rect 24032 20927 24084 20936
rect 24032 20893 24041 20927
rect 24041 20893 24075 20927
rect 24075 20893 24084 20927
rect 24032 20884 24084 20893
rect 24400 20884 24452 20936
rect 23388 20816 23440 20868
rect 21640 20748 21692 20800
rect 22192 20748 22244 20800
rect 22560 20748 22612 20800
rect 23664 20748 23716 20800
rect 23940 20748 23992 20800
rect 4922 20646 4974 20698
rect 4986 20646 5038 20698
rect 5050 20646 5102 20698
rect 5114 20646 5166 20698
rect 5178 20646 5230 20698
rect 5242 20646 5294 20698
rect 10922 20646 10974 20698
rect 10986 20646 11038 20698
rect 11050 20646 11102 20698
rect 11114 20646 11166 20698
rect 11178 20646 11230 20698
rect 11242 20646 11294 20698
rect 16922 20646 16974 20698
rect 16986 20646 17038 20698
rect 17050 20646 17102 20698
rect 17114 20646 17166 20698
rect 17178 20646 17230 20698
rect 17242 20646 17294 20698
rect 22922 20646 22974 20698
rect 22986 20646 23038 20698
rect 23050 20646 23102 20698
rect 23114 20646 23166 20698
rect 23178 20646 23230 20698
rect 23242 20646 23294 20698
rect 28922 20646 28974 20698
rect 28986 20646 29038 20698
rect 29050 20646 29102 20698
rect 29114 20646 29166 20698
rect 29178 20646 29230 20698
rect 29242 20646 29294 20698
rect 4160 20587 4212 20596
rect 4160 20553 4169 20587
rect 4169 20553 4203 20587
rect 4203 20553 4212 20587
rect 4160 20544 4212 20553
rect 5356 20544 5408 20596
rect 6644 20544 6696 20596
rect 6920 20544 6972 20596
rect 7472 20587 7524 20596
rect 7472 20553 7481 20587
rect 7481 20553 7515 20587
rect 7515 20553 7524 20587
rect 7472 20544 7524 20553
rect 5540 20408 5592 20460
rect 6092 20408 6144 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 8484 20451 8536 20460
rect 8484 20417 8518 20451
rect 8518 20417 8536 20451
rect 8484 20408 8536 20417
rect 8760 20408 8812 20460
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 6828 20340 6880 20392
rect 10784 20408 10836 20460
rect 1860 20272 1912 20324
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 11704 20408 11756 20460
rect 12440 20476 12492 20528
rect 12624 20544 12676 20596
rect 14096 20544 14148 20596
rect 16028 20544 16080 20596
rect 16120 20544 16172 20596
rect 18052 20544 18104 20596
rect 12164 20451 12216 20460
rect 12164 20417 12198 20451
rect 12198 20417 12216 20451
rect 12164 20408 12216 20417
rect 16672 20476 16724 20528
rect 17592 20476 17644 20528
rect 13728 20408 13780 20460
rect 13636 20340 13688 20392
rect 14648 20408 14700 20460
rect 14740 20408 14792 20460
rect 14832 20408 14884 20460
rect 15568 20408 15620 20460
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 6368 20247 6420 20256
rect 6368 20213 6377 20247
rect 6377 20213 6411 20247
rect 6411 20213 6420 20247
rect 6368 20204 6420 20213
rect 14004 20272 14056 20324
rect 16028 20408 16080 20460
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 17868 20408 17920 20460
rect 18604 20476 18656 20528
rect 19248 20476 19300 20528
rect 20720 20519 20772 20528
rect 20720 20485 20729 20519
rect 20729 20485 20763 20519
rect 20763 20485 20772 20519
rect 20720 20476 20772 20485
rect 20996 20476 21048 20528
rect 21548 20544 21600 20596
rect 21732 20544 21784 20596
rect 21824 20544 21876 20596
rect 22192 20544 22244 20596
rect 23296 20544 23348 20596
rect 24124 20544 24176 20596
rect 21364 20408 21416 20460
rect 16488 20340 16540 20392
rect 15844 20247 15896 20256
rect 15844 20213 15853 20247
rect 15853 20213 15887 20247
rect 15887 20213 15896 20247
rect 15844 20204 15896 20213
rect 16028 20204 16080 20256
rect 17500 20204 17552 20256
rect 17776 20204 17828 20256
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 19708 20204 19760 20256
rect 20904 20340 20956 20392
rect 21732 20340 21784 20392
rect 20812 20272 20864 20324
rect 21916 20408 21968 20460
rect 22100 20340 22152 20392
rect 22560 20451 22612 20460
rect 22560 20417 22569 20451
rect 22569 20417 22603 20451
rect 22603 20417 22612 20451
rect 22560 20408 22612 20417
rect 23480 20408 23532 20460
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 24032 20408 24084 20460
rect 24676 20451 24728 20460
rect 24676 20417 24685 20451
rect 24685 20417 24719 20451
rect 24719 20417 24728 20451
rect 24676 20408 24728 20417
rect 23112 20340 23164 20392
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23296 20340 23348 20349
rect 24400 20340 24452 20392
rect 23572 20272 23624 20324
rect 22468 20204 22520 20256
rect 22928 20204 22980 20256
rect 23756 20204 23808 20256
rect 4182 20102 4234 20154
rect 4246 20102 4298 20154
rect 4310 20102 4362 20154
rect 4374 20102 4426 20154
rect 4438 20102 4490 20154
rect 4502 20102 4554 20154
rect 10182 20102 10234 20154
rect 10246 20102 10298 20154
rect 10310 20102 10362 20154
rect 10374 20102 10426 20154
rect 10438 20102 10490 20154
rect 10502 20102 10554 20154
rect 16182 20102 16234 20154
rect 16246 20102 16298 20154
rect 16310 20102 16362 20154
rect 16374 20102 16426 20154
rect 16438 20102 16490 20154
rect 16502 20102 16554 20154
rect 22182 20102 22234 20154
rect 22246 20102 22298 20154
rect 22310 20102 22362 20154
rect 22374 20102 22426 20154
rect 22438 20102 22490 20154
rect 22502 20102 22554 20154
rect 28182 20102 28234 20154
rect 28246 20102 28298 20154
rect 28310 20102 28362 20154
rect 28374 20102 28426 20154
rect 28438 20102 28490 20154
rect 28502 20102 28554 20154
rect 5540 20043 5592 20052
rect 5540 20009 5549 20043
rect 5549 20009 5583 20043
rect 5583 20009 5592 20043
rect 5540 20000 5592 20009
rect 6368 20000 6420 20052
rect 6828 20000 6880 20052
rect 10784 19932 10836 19984
rect 11428 20043 11480 20052
rect 11428 20009 11437 20043
rect 11437 20009 11471 20043
rect 11471 20009 11480 20043
rect 11428 20000 11480 20009
rect 12716 20000 12768 20052
rect 16672 20000 16724 20052
rect 8300 19796 8352 19848
rect 9956 19796 10008 19848
rect 10600 19796 10652 19848
rect 10876 19839 10928 19848
rect 10876 19805 10885 19839
rect 10885 19805 10919 19839
rect 10919 19805 10928 19839
rect 10876 19796 10928 19805
rect 12716 19864 12768 19916
rect 15292 19864 15344 19916
rect 15752 19932 15804 19984
rect 19064 19975 19116 19984
rect 19064 19941 19073 19975
rect 19073 19941 19107 19975
rect 19107 19941 19116 19975
rect 19064 19932 19116 19941
rect 19156 19932 19208 19984
rect 19340 19932 19392 19984
rect 22100 20000 22152 20052
rect 14004 19796 14056 19848
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 20904 19864 20956 19916
rect 21824 19932 21876 19984
rect 1676 19660 1728 19712
rect 11980 19660 12032 19712
rect 16028 19660 16080 19712
rect 16764 19796 16816 19848
rect 17408 19796 17460 19848
rect 18604 19796 18656 19848
rect 19340 19796 19392 19848
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19892 19796 19944 19848
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 20996 19796 21048 19848
rect 21456 19864 21508 19916
rect 21732 19796 21784 19848
rect 22652 20000 22704 20052
rect 22928 19932 22980 19984
rect 24400 19932 24452 19984
rect 24492 19932 24544 19984
rect 17500 19728 17552 19780
rect 20260 19728 20312 19780
rect 18880 19703 18932 19712
rect 18880 19669 18915 19703
rect 18915 19669 18932 19703
rect 18880 19660 18932 19669
rect 19248 19660 19300 19712
rect 20444 19771 20496 19780
rect 20444 19737 20453 19771
rect 20453 19737 20487 19771
rect 20487 19737 20496 19771
rect 20444 19728 20496 19737
rect 20720 19728 20772 19780
rect 21272 19728 21324 19780
rect 21548 19728 21600 19780
rect 21640 19728 21692 19780
rect 22652 19796 22704 19848
rect 23112 19839 23164 19848
rect 23112 19805 23121 19839
rect 23121 19805 23155 19839
rect 23155 19805 23164 19839
rect 23112 19796 23164 19805
rect 23664 19796 23716 19848
rect 23388 19728 23440 19780
rect 24032 19796 24084 19848
rect 24492 19796 24544 19848
rect 21088 19660 21140 19712
rect 21456 19703 21508 19712
rect 21456 19669 21465 19703
rect 21465 19669 21499 19703
rect 21499 19669 21508 19703
rect 21456 19660 21508 19669
rect 21824 19703 21876 19712
rect 21824 19669 21833 19703
rect 21833 19669 21867 19703
rect 21867 19669 21876 19703
rect 21824 19660 21876 19669
rect 21916 19660 21968 19712
rect 23480 19660 23532 19712
rect 26700 19839 26752 19848
rect 26700 19805 26709 19839
rect 26709 19805 26743 19839
rect 26743 19805 26752 19839
rect 26700 19796 26752 19805
rect 24768 19660 24820 19712
rect 26608 19703 26660 19712
rect 26608 19669 26617 19703
rect 26617 19669 26651 19703
rect 26651 19669 26660 19703
rect 26608 19660 26660 19669
rect 4922 19558 4974 19610
rect 4986 19558 5038 19610
rect 5050 19558 5102 19610
rect 5114 19558 5166 19610
rect 5178 19558 5230 19610
rect 5242 19558 5294 19610
rect 10922 19558 10974 19610
rect 10986 19558 11038 19610
rect 11050 19558 11102 19610
rect 11114 19558 11166 19610
rect 11178 19558 11230 19610
rect 11242 19558 11294 19610
rect 16922 19558 16974 19610
rect 16986 19558 17038 19610
rect 17050 19558 17102 19610
rect 17114 19558 17166 19610
rect 17178 19558 17230 19610
rect 17242 19558 17294 19610
rect 22922 19558 22974 19610
rect 22986 19558 23038 19610
rect 23050 19558 23102 19610
rect 23114 19558 23166 19610
rect 23178 19558 23230 19610
rect 23242 19558 23294 19610
rect 28922 19558 28974 19610
rect 28986 19558 29038 19610
rect 29050 19558 29102 19610
rect 29114 19558 29166 19610
rect 29178 19558 29230 19610
rect 29242 19558 29294 19610
rect 7564 19456 7616 19508
rect 14188 19456 14240 19508
rect 15292 19456 15344 19508
rect 14832 19388 14884 19440
rect 15752 19388 15804 19440
rect 15844 19388 15896 19440
rect 16488 19456 16540 19508
rect 19156 19456 19208 19508
rect 22560 19456 22612 19508
rect 23756 19456 23808 19508
rect 19248 19388 19300 19440
rect 21456 19388 21508 19440
rect 3332 19320 3384 19372
rect 15568 19320 15620 19372
rect 17408 19320 17460 19372
rect 17684 19363 17736 19372
rect 17684 19329 17693 19363
rect 17693 19329 17727 19363
rect 17727 19329 17736 19363
rect 17684 19320 17736 19329
rect 26608 19388 26660 19440
rect 4620 19252 4672 19304
rect 5080 19252 5132 19304
rect 15200 19184 15252 19236
rect 16580 19252 16632 19304
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 3792 19159 3844 19168
rect 3792 19125 3801 19159
rect 3801 19125 3835 19159
rect 3835 19125 3844 19159
rect 3792 19116 3844 19125
rect 4068 19116 4120 19168
rect 4712 19116 4764 19168
rect 10048 19116 10100 19168
rect 15476 19116 15528 19168
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 17316 19184 17368 19236
rect 18236 19184 18288 19236
rect 18604 19184 18656 19236
rect 20444 19320 20496 19372
rect 20904 19320 20956 19372
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 22100 19320 22152 19372
rect 22652 19320 22704 19372
rect 24952 19363 25004 19372
rect 24952 19329 24961 19363
rect 24961 19329 24995 19363
rect 24995 19329 25004 19363
rect 24952 19320 25004 19329
rect 25044 19363 25096 19372
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 29644 19320 29696 19372
rect 20628 19295 20680 19304
rect 20628 19261 20637 19295
rect 20637 19261 20671 19295
rect 20671 19261 20680 19295
rect 20628 19252 20680 19261
rect 21180 19252 21232 19304
rect 21272 19252 21324 19304
rect 21916 19252 21968 19304
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 17592 19116 17644 19168
rect 18880 19116 18932 19168
rect 21548 19116 21600 19168
rect 23480 19116 23532 19168
rect 24400 19116 24452 19168
rect 30932 19116 30984 19168
rect 4182 19014 4234 19066
rect 4246 19014 4298 19066
rect 4310 19014 4362 19066
rect 4374 19014 4426 19066
rect 4438 19014 4490 19066
rect 4502 19014 4554 19066
rect 10182 19014 10234 19066
rect 10246 19014 10298 19066
rect 10310 19014 10362 19066
rect 10374 19014 10426 19066
rect 10438 19014 10490 19066
rect 10502 19014 10554 19066
rect 16182 19014 16234 19066
rect 16246 19014 16298 19066
rect 16310 19014 16362 19066
rect 16374 19014 16426 19066
rect 16438 19014 16490 19066
rect 16502 19014 16554 19066
rect 22182 19014 22234 19066
rect 22246 19014 22298 19066
rect 22310 19014 22362 19066
rect 22374 19014 22426 19066
rect 22438 19014 22490 19066
rect 22502 19014 22554 19066
rect 28182 19014 28234 19066
rect 28246 19014 28298 19066
rect 28310 19014 28362 19066
rect 28374 19014 28426 19066
rect 28438 19014 28490 19066
rect 28502 19014 28554 19066
rect 3332 18912 3384 18964
rect 4528 18912 4580 18964
rect 4712 18844 4764 18896
rect 6552 18912 6604 18964
rect 16304 18912 16356 18964
rect 3976 18776 4028 18828
rect 5080 18776 5132 18828
rect 15108 18844 15160 18896
rect 19800 18912 19852 18964
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 4804 18708 4856 18760
rect 2596 18640 2648 18692
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 6460 18572 6512 18624
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 9772 18708 9824 18760
rect 6828 18640 6880 18692
rect 14096 18708 14148 18760
rect 14188 18708 14240 18760
rect 14740 18751 14792 18760
rect 14740 18717 14749 18751
rect 14749 18717 14783 18751
rect 14783 18717 14792 18751
rect 14740 18708 14792 18717
rect 15660 18776 15712 18828
rect 16488 18819 16540 18828
rect 16488 18785 16497 18819
rect 16497 18785 16531 18819
rect 16531 18785 16540 18819
rect 16488 18776 16540 18785
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 17408 18776 17460 18828
rect 17500 18776 17552 18828
rect 17960 18776 18012 18828
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 17408 18640 17460 18692
rect 17868 18708 17920 18760
rect 19708 18708 19760 18760
rect 21732 18912 21784 18964
rect 24492 18955 24544 18964
rect 24492 18921 24501 18955
rect 24501 18921 24535 18955
rect 24535 18921 24544 18955
rect 24492 18912 24544 18921
rect 25320 18955 25372 18964
rect 25320 18921 25329 18955
rect 25329 18921 25363 18955
rect 25363 18921 25372 18955
rect 25320 18912 25372 18921
rect 21824 18844 21876 18896
rect 21640 18819 21692 18828
rect 21640 18785 21649 18819
rect 21649 18785 21683 18819
rect 21683 18785 21692 18819
rect 21640 18776 21692 18785
rect 23572 18844 23624 18896
rect 24676 18844 24728 18896
rect 21548 18708 21600 18760
rect 25136 18751 25188 18760
rect 25136 18717 25145 18751
rect 25145 18717 25179 18751
rect 25179 18717 25188 18751
rect 25136 18708 25188 18717
rect 21272 18683 21324 18692
rect 21272 18649 21281 18683
rect 21281 18649 21315 18683
rect 21315 18649 21324 18683
rect 21272 18640 21324 18649
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 17684 18572 17736 18624
rect 21824 18615 21876 18624
rect 21824 18581 21833 18615
rect 21833 18581 21867 18615
rect 21867 18581 21876 18615
rect 21824 18572 21876 18581
rect 24676 18572 24728 18624
rect 24860 18572 24912 18624
rect 4922 18470 4974 18522
rect 4986 18470 5038 18522
rect 5050 18470 5102 18522
rect 5114 18470 5166 18522
rect 5178 18470 5230 18522
rect 5242 18470 5294 18522
rect 10922 18470 10974 18522
rect 10986 18470 11038 18522
rect 11050 18470 11102 18522
rect 11114 18470 11166 18522
rect 11178 18470 11230 18522
rect 11242 18470 11294 18522
rect 16922 18470 16974 18522
rect 16986 18470 17038 18522
rect 17050 18470 17102 18522
rect 17114 18470 17166 18522
rect 17178 18470 17230 18522
rect 17242 18470 17294 18522
rect 22922 18470 22974 18522
rect 22986 18470 23038 18522
rect 23050 18470 23102 18522
rect 23114 18470 23166 18522
rect 23178 18470 23230 18522
rect 23242 18470 23294 18522
rect 28922 18470 28974 18522
rect 28986 18470 29038 18522
rect 29050 18470 29102 18522
rect 29114 18470 29166 18522
rect 29178 18470 29230 18522
rect 29242 18470 29294 18522
rect 2228 18368 2280 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 3792 18368 3844 18420
rect 4252 18368 4304 18420
rect 4620 18368 4672 18420
rect 4712 18368 4764 18420
rect 2412 18275 2464 18284
rect 2412 18241 2446 18275
rect 2446 18241 2464 18275
rect 2412 18232 2464 18241
rect 4528 18300 4580 18352
rect 5448 18232 5500 18284
rect 6552 18368 6604 18420
rect 6736 18368 6788 18420
rect 3240 18164 3292 18216
rect 6828 18164 6880 18216
rect 3056 18028 3108 18080
rect 6460 18096 6512 18148
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 4068 18028 4120 18080
rect 5908 18071 5960 18080
rect 5908 18037 5917 18071
rect 5917 18037 5951 18071
rect 5951 18037 5960 18071
rect 5908 18028 5960 18037
rect 8392 18343 8444 18352
rect 8392 18309 8401 18343
rect 8401 18309 8435 18343
rect 8435 18309 8444 18343
rect 8392 18300 8444 18309
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 9128 18368 9180 18420
rect 15936 18368 15988 18420
rect 16672 18368 16724 18420
rect 12716 18343 12768 18352
rect 12716 18309 12739 18343
rect 12739 18309 12768 18343
rect 12716 18300 12768 18309
rect 15844 18300 15896 18352
rect 8116 18164 8168 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 11612 18232 11664 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 15200 18232 15252 18284
rect 16028 18232 16080 18284
rect 16488 18300 16540 18352
rect 16764 18300 16816 18352
rect 18420 18300 18472 18352
rect 23388 18300 23440 18352
rect 23480 18343 23532 18352
rect 23480 18309 23489 18343
rect 23489 18309 23523 18343
rect 23523 18309 23532 18343
rect 23480 18300 23532 18309
rect 23572 18300 23624 18352
rect 16304 18232 16356 18284
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 18972 18232 19024 18284
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 10600 18164 10652 18216
rect 14280 18207 14332 18216
rect 14280 18173 14289 18207
rect 14289 18173 14323 18207
rect 14323 18173 14332 18207
rect 14280 18164 14332 18173
rect 15476 18164 15528 18216
rect 15936 18164 15988 18216
rect 16580 18164 16632 18216
rect 17500 18164 17552 18216
rect 9956 18096 10008 18148
rect 17776 18164 17828 18216
rect 19708 18232 19760 18284
rect 21548 18232 21600 18284
rect 20720 18164 20772 18216
rect 24400 18343 24452 18352
rect 24400 18309 24409 18343
rect 24409 18309 24443 18343
rect 24443 18309 24452 18343
rect 24400 18300 24452 18309
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 24952 18232 25004 18284
rect 14556 18028 14608 18080
rect 15108 18028 15160 18080
rect 19616 18096 19668 18148
rect 26700 18164 26752 18216
rect 26976 18164 27028 18216
rect 24860 18139 24912 18148
rect 24860 18105 24884 18139
rect 24884 18105 24912 18139
rect 24860 18096 24912 18105
rect 20076 18028 20128 18080
rect 21272 18028 21324 18080
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 23112 18071 23164 18080
rect 23112 18037 23121 18071
rect 23121 18037 23155 18071
rect 23155 18037 23164 18071
rect 23112 18028 23164 18037
rect 24032 18071 24084 18080
rect 24032 18037 24041 18071
rect 24041 18037 24075 18071
rect 24075 18037 24084 18071
rect 24032 18028 24084 18037
rect 24676 18028 24728 18080
rect 26332 18028 26384 18080
rect 27068 18028 27120 18080
rect 27620 18028 27672 18080
rect 4182 17926 4234 17978
rect 4246 17926 4298 17978
rect 4310 17926 4362 17978
rect 4374 17926 4426 17978
rect 4438 17926 4490 17978
rect 4502 17926 4554 17978
rect 10182 17926 10234 17978
rect 10246 17926 10298 17978
rect 10310 17926 10362 17978
rect 10374 17926 10426 17978
rect 10438 17926 10490 17978
rect 10502 17926 10554 17978
rect 16182 17926 16234 17978
rect 16246 17926 16298 17978
rect 16310 17926 16362 17978
rect 16374 17926 16426 17978
rect 16438 17926 16490 17978
rect 16502 17926 16554 17978
rect 22182 17926 22234 17978
rect 22246 17926 22298 17978
rect 22310 17926 22362 17978
rect 22374 17926 22426 17978
rect 22438 17926 22490 17978
rect 22502 17926 22554 17978
rect 28182 17926 28234 17978
rect 28246 17926 28298 17978
rect 28310 17926 28362 17978
rect 28374 17926 28426 17978
rect 28438 17926 28490 17978
rect 28502 17926 28554 17978
rect 2412 17824 2464 17876
rect 5448 17824 5500 17876
rect 4804 17688 4856 17740
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 8208 17756 8260 17808
rect 12256 17824 12308 17876
rect 9680 17756 9732 17808
rect 3608 17620 3660 17672
rect 9588 17688 9640 17740
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 17224 17824 17276 17876
rect 15200 17756 15252 17808
rect 15936 17756 15988 17808
rect 9956 17620 10008 17672
rect 11888 17688 11940 17740
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13636 17688 13688 17740
rect 14556 17731 14608 17740
rect 14556 17697 14565 17731
rect 14565 17697 14599 17731
rect 14599 17697 14608 17731
rect 14556 17688 14608 17697
rect 14740 17731 14792 17740
rect 14740 17697 14749 17731
rect 14749 17697 14783 17731
rect 14783 17697 14792 17731
rect 14740 17688 14792 17697
rect 15476 17688 15528 17740
rect 15660 17688 15712 17740
rect 5908 17552 5960 17604
rect 6552 17552 6604 17604
rect 11612 17620 11664 17672
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 16856 17756 16908 17808
rect 16764 17731 16816 17740
rect 16764 17697 16773 17731
rect 16773 17697 16807 17731
rect 16807 17697 16816 17731
rect 16764 17688 16816 17697
rect 17500 17688 17552 17740
rect 8116 17484 8168 17536
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 10140 17484 10192 17536
rect 10416 17527 10468 17536
rect 10416 17493 10425 17527
rect 10425 17493 10459 17527
rect 10459 17493 10468 17527
rect 10416 17484 10468 17493
rect 11336 17484 11388 17536
rect 11612 17484 11664 17536
rect 14096 17552 14148 17604
rect 14372 17484 14424 17536
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14464 17484 14516 17493
rect 15568 17552 15620 17604
rect 15752 17552 15804 17604
rect 15936 17552 15988 17604
rect 17960 17663 18012 17672
rect 17960 17629 17969 17663
rect 17969 17629 18003 17663
rect 18003 17629 18012 17663
rect 17960 17620 18012 17629
rect 19248 17824 19300 17876
rect 19892 17824 19944 17876
rect 25136 17824 25188 17876
rect 26332 17824 26384 17876
rect 18696 17688 18748 17740
rect 18236 17552 18288 17604
rect 19340 17688 19392 17740
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 19156 17620 19208 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 19892 17620 19944 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 23388 17731 23440 17740
rect 23388 17697 23397 17731
rect 23397 17697 23431 17731
rect 23431 17697 23440 17731
rect 23388 17688 23440 17697
rect 25044 17688 25096 17740
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 21824 17620 21876 17672
rect 22100 17620 22152 17672
rect 17868 17484 17920 17536
rect 18972 17484 19024 17536
rect 20260 17595 20312 17604
rect 20260 17561 20269 17595
rect 20269 17561 20303 17595
rect 20303 17561 20312 17595
rect 20260 17552 20312 17561
rect 21732 17595 21784 17604
rect 21732 17561 21741 17595
rect 21741 17561 21775 17595
rect 21775 17561 21784 17595
rect 21732 17552 21784 17561
rect 22284 17552 22336 17604
rect 24768 17620 24820 17672
rect 25504 17663 25556 17672
rect 25504 17629 25513 17663
rect 25513 17629 25547 17663
rect 25547 17629 25556 17663
rect 25504 17620 25556 17629
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 21088 17484 21140 17536
rect 22560 17484 22612 17536
rect 23112 17552 23164 17604
rect 23572 17595 23624 17604
rect 23572 17561 23581 17595
rect 23581 17561 23615 17595
rect 23615 17561 23624 17595
rect 23572 17552 23624 17561
rect 27068 17552 27120 17604
rect 4922 17382 4974 17434
rect 4986 17382 5038 17434
rect 5050 17382 5102 17434
rect 5114 17382 5166 17434
rect 5178 17382 5230 17434
rect 5242 17382 5294 17434
rect 10922 17382 10974 17434
rect 10986 17382 11038 17434
rect 11050 17382 11102 17434
rect 11114 17382 11166 17434
rect 11178 17382 11230 17434
rect 11242 17382 11294 17434
rect 16922 17382 16974 17434
rect 16986 17382 17038 17434
rect 17050 17382 17102 17434
rect 17114 17382 17166 17434
rect 17178 17382 17230 17434
rect 17242 17382 17294 17434
rect 22922 17382 22974 17434
rect 22986 17382 23038 17434
rect 23050 17382 23102 17434
rect 23114 17382 23166 17434
rect 23178 17382 23230 17434
rect 23242 17382 23294 17434
rect 28922 17382 28974 17434
rect 28986 17382 29038 17434
rect 29050 17382 29102 17434
rect 29114 17382 29166 17434
rect 29178 17382 29230 17434
rect 29242 17382 29294 17434
rect 6552 17280 6604 17332
rect 6736 17280 6788 17332
rect 8300 17280 8352 17332
rect 8392 17280 8444 17332
rect 8116 17212 8168 17264
rect 6460 17076 6512 17128
rect 6828 17076 6880 17128
rect 8208 17187 8260 17196
rect 8208 17153 8217 17187
rect 8217 17153 8251 17187
rect 8251 17153 8260 17187
rect 8208 17144 8260 17153
rect 8484 17144 8536 17196
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 9128 17212 9180 17264
rect 9588 17212 9640 17264
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 10416 17280 10468 17332
rect 11612 17280 11664 17332
rect 10600 17255 10652 17264
rect 10600 17221 10609 17255
rect 10609 17221 10643 17255
rect 10643 17221 10652 17255
rect 10600 17212 10652 17221
rect 12164 17280 12216 17332
rect 15200 17323 15252 17332
rect 15200 17289 15209 17323
rect 15209 17289 15243 17323
rect 15243 17289 15252 17323
rect 15200 17280 15252 17289
rect 16672 17280 16724 17332
rect 18420 17323 18472 17332
rect 18420 17289 18429 17323
rect 18429 17289 18463 17323
rect 18463 17289 18472 17323
rect 18420 17280 18472 17289
rect 19524 17323 19576 17332
rect 19524 17289 19533 17323
rect 19533 17289 19567 17323
rect 19567 17289 19576 17323
rect 19524 17280 19576 17289
rect 20260 17280 20312 17332
rect 15108 17212 15160 17264
rect 16764 17212 16816 17264
rect 17684 17255 17736 17264
rect 17684 17221 17693 17255
rect 17693 17221 17727 17255
rect 17727 17221 17736 17255
rect 17684 17212 17736 17221
rect 19064 17212 19116 17264
rect 24032 17280 24084 17332
rect 21364 17212 21416 17264
rect 22652 17212 22704 17264
rect 23480 17212 23532 17264
rect 24768 17280 24820 17332
rect 25504 17280 25556 17332
rect 10048 17076 10100 17128
rect 11428 17144 11480 17196
rect 11520 17187 11572 17196
rect 11520 17153 11529 17187
rect 11529 17153 11563 17187
rect 11563 17153 11572 17187
rect 11520 17144 11572 17153
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11152 17076 11204 17128
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 16488 17187 16540 17196
rect 16488 17153 16497 17187
rect 16497 17153 16531 17187
rect 16531 17153 16540 17187
rect 16488 17144 16540 17153
rect 13452 17119 13504 17128
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 13636 17119 13688 17128
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 16580 17076 16632 17128
rect 17868 17144 17920 17196
rect 18144 17144 18196 17196
rect 17408 17008 17460 17060
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 22100 17144 22152 17196
rect 22560 17144 22612 17196
rect 22928 17144 22980 17196
rect 23664 17144 23716 17196
rect 26976 17144 27028 17196
rect 18420 17076 18472 17128
rect 18972 17076 19024 17128
rect 19064 17119 19116 17128
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 20904 17076 20956 17128
rect 12256 16940 12308 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 16764 16940 16816 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 20720 16940 20772 16992
rect 20996 17008 21048 17060
rect 21272 17119 21324 17128
rect 21272 17085 21281 17119
rect 21281 17085 21315 17119
rect 21315 17085 21324 17119
rect 21272 17076 21324 17085
rect 22284 17008 22336 17060
rect 23020 17076 23072 17128
rect 23388 17076 23440 17128
rect 23572 17008 23624 17060
rect 23940 17119 23992 17128
rect 23940 17085 23949 17119
rect 23949 17085 23983 17119
rect 23983 17085 23992 17119
rect 23940 17076 23992 17085
rect 24860 17008 24912 17060
rect 22008 16983 22060 16992
rect 22008 16949 22032 16983
rect 22032 16949 22060 16983
rect 22008 16940 22060 16949
rect 22652 16940 22704 16992
rect 25504 16983 25556 16992
rect 25504 16949 25513 16983
rect 25513 16949 25547 16983
rect 25547 16949 25556 16983
rect 25504 16940 25556 16949
rect 27160 16940 27212 16992
rect 4182 16838 4234 16890
rect 4246 16838 4298 16890
rect 4310 16838 4362 16890
rect 4374 16838 4426 16890
rect 4438 16838 4490 16890
rect 4502 16838 4554 16890
rect 10182 16838 10234 16890
rect 10246 16838 10298 16890
rect 10310 16838 10362 16890
rect 10374 16838 10426 16890
rect 10438 16838 10490 16890
rect 10502 16838 10554 16890
rect 16182 16838 16234 16890
rect 16246 16838 16298 16890
rect 16310 16838 16362 16890
rect 16374 16838 16426 16890
rect 16438 16838 16490 16890
rect 16502 16838 16554 16890
rect 22182 16838 22234 16890
rect 22246 16838 22298 16890
rect 22310 16838 22362 16890
rect 22374 16838 22426 16890
rect 22438 16838 22490 16890
rect 22502 16838 22554 16890
rect 28182 16838 28234 16890
rect 28246 16838 28298 16890
rect 28310 16838 28362 16890
rect 28374 16838 28426 16890
rect 28438 16838 28490 16890
rect 28502 16838 28554 16890
rect 3884 16736 3936 16788
rect 8024 16736 8076 16788
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 11152 16779 11204 16788
rect 11152 16745 11161 16779
rect 11161 16745 11195 16779
rect 11195 16745 11204 16779
rect 11152 16736 11204 16745
rect 6828 16668 6880 16720
rect 14096 16736 14148 16788
rect 14372 16736 14424 16788
rect 15936 16736 15988 16788
rect 16672 16736 16724 16788
rect 18052 16736 18104 16788
rect 19064 16736 19116 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 20720 16736 20772 16788
rect 21732 16736 21784 16788
rect 22376 16736 22428 16788
rect 23020 16736 23072 16788
rect 23112 16736 23164 16788
rect 11520 16668 11572 16720
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 4620 16600 4672 16652
rect 9588 16600 9640 16652
rect 2320 16439 2372 16448
rect 2320 16405 2329 16439
rect 2329 16405 2363 16439
rect 2363 16405 2372 16439
rect 2320 16396 2372 16405
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 11428 16600 11480 16652
rect 11888 16600 11940 16652
rect 11704 16532 11756 16584
rect 10784 16507 10836 16516
rect 10784 16473 10793 16507
rect 10793 16473 10827 16507
rect 10827 16473 10836 16507
rect 10784 16464 10836 16473
rect 11152 16396 11204 16448
rect 11336 16396 11388 16448
rect 11888 16396 11940 16448
rect 15292 16600 15344 16652
rect 14188 16464 14240 16516
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 14740 16532 14792 16584
rect 15200 16396 15252 16448
rect 15660 16507 15712 16516
rect 15660 16473 15669 16507
rect 15669 16473 15703 16507
rect 15703 16473 15712 16507
rect 15660 16464 15712 16473
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 17592 16668 17644 16720
rect 18420 16643 18472 16652
rect 15752 16396 15804 16448
rect 18420 16609 18429 16643
rect 18429 16609 18463 16643
rect 18463 16609 18472 16643
rect 18420 16600 18472 16609
rect 18696 16532 18748 16584
rect 19248 16600 19300 16652
rect 23204 16668 23256 16720
rect 23940 16736 23992 16788
rect 25504 16736 25556 16788
rect 27620 16779 27672 16788
rect 27620 16745 27629 16779
rect 27629 16745 27663 16779
rect 27663 16745 27672 16779
rect 27620 16736 27672 16745
rect 23572 16668 23624 16720
rect 19248 16507 19300 16516
rect 19248 16473 19257 16507
rect 19257 16473 19291 16507
rect 19291 16473 19300 16507
rect 19248 16464 19300 16473
rect 20076 16464 20128 16516
rect 24400 16643 24452 16652
rect 24400 16609 24409 16643
rect 24409 16609 24443 16643
rect 24443 16609 24452 16643
rect 24400 16600 24452 16609
rect 26240 16600 26292 16652
rect 22100 16532 22152 16584
rect 22928 16575 22980 16584
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 23112 16532 23164 16584
rect 23204 16575 23256 16584
rect 23204 16541 23213 16575
rect 23213 16541 23247 16575
rect 23247 16541 23256 16575
rect 23204 16532 23256 16541
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 19156 16396 19208 16448
rect 19340 16396 19392 16448
rect 19892 16396 19944 16448
rect 21364 16464 21416 16516
rect 24032 16532 24084 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 27160 16532 27212 16584
rect 20996 16396 21048 16448
rect 24308 16464 24360 16516
rect 26516 16396 26568 16448
rect 4922 16294 4974 16346
rect 4986 16294 5038 16346
rect 5050 16294 5102 16346
rect 5114 16294 5166 16346
rect 5178 16294 5230 16346
rect 5242 16294 5294 16346
rect 10922 16294 10974 16346
rect 10986 16294 11038 16346
rect 11050 16294 11102 16346
rect 11114 16294 11166 16346
rect 11178 16294 11230 16346
rect 11242 16294 11294 16346
rect 16922 16294 16974 16346
rect 16986 16294 17038 16346
rect 17050 16294 17102 16346
rect 17114 16294 17166 16346
rect 17178 16294 17230 16346
rect 17242 16294 17294 16346
rect 22922 16294 22974 16346
rect 22986 16294 23038 16346
rect 23050 16294 23102 16346
rect 23114 16294 23166 16346
rect 23178 16294 23230 16346
rect 23242 16294 23294 16346
rect 28922 16294 28974 16346
rect 28986 16294 29038 16346
rect 29050 16294 29102 16346
rect 29114 16294 29166 16346
rect 29178 16294 29230 16346
rect 29242 16294 29294 16346
rect 4344 16192 4396 16244
rect 6644 16192 6696 16244
rect 8392 16192 8444 16244
rect 2320 16124 2372 16176
rect 3884 16167 3936 16176
rect 3884 16133 3893 16167
rect 3893 16133 3927 16167
rect 3927 16133 3936 16167
rect 3884 16124 3936 16133
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 4712 16124 4764 16176
rect 3976 16031 4028 16040
rect 3976 15997 3985 16031
rect 3985 15997 4019 16031
rect 4019 15997 4028 16031
rect 3976 15988 4028 15997
rect 5448 16056 5500 16108
rect 10324 16192 10376 16244
rect 11336 16192 11388 16244
rect 15660 16192 15712 16244
rect 16764 16192 16816 16244
rect 18144 16192 18196 16244
rect 10968 16124 11020 16176
rect 1860 15895 1912 15904
rect 1860 15861 1869 15895
rect 1869 15861 1903 15895
rect 1903 15861 1912 15895
rect 1860 15852 1912 15861
rect 3240 15852 3292 15904
rect 6828 15988 6880 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 7932 15988 7984 16040
rect 9772 15988 9824 16040
rect 11428 15988 11480 16040
rect 7288 15920 7340 15972
rect 12624 16056 12676 16108
rect 16028 16124 16080 16176
rect 18328 16192 18380 16244
rect 18512 16192 18564 16244
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 14740 15920 14792 15972
rect 4804 15852 4856 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 14832 15852 14884 15904
rect 15108 15852 15160 15904
rect 18236 16056 18288 16108
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 18788 16192 18840 16244
rect 19156 16056 19208 16108
rect 19616 16056 19668 16108
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 21364 16235 21416 16244
rect 21364 16201 21373 16235
rect 21373 16201 21407 16235
rect 21407 16201 21416 16235
rect 21364 16192 21416 16201
rect 23572 16192 23624 16244
rect 24860 16192 24912 16244
rect 22100 16124 22152 16176
rect 20904 16056 20956 16108
rect 22008 16056 22060 16108
rect 25504 16124 25556 16176
rect 23848 16099 23900 16108
rect 23848 16065 23857 16099
rect 23857 16065 23891 16099
rect 23891 16065 23900 16099
rect 23848 16056 23900 16065
rect 24400 16056 24452 16108
rect 26148 16099 26200 16108
rect 26148 16065 26157 16099
rect 26157 16065 26191 16099
rect 26191 16065 26200 16099
rect 26148 16056 26200 16065
rect 18696 15920 18748 15972
rect 19616 15920 19668 15972
rect 22376 15988 22428 16040
rect 26516 16099 26568 16108
rect 26516 16065 26525 16099
rect 26525 16065 26559 16099
rect 26559 16065 26568 16099
rect 26516 16056 26568 16065
rect 27068 16056 27120 16108
rect 23388 15920 23440 15972
rect 27528 15988 27580 16040
rect 25688 15852 25740 15904
rect 26700 15895 26752 15904
rect 26700 15861 26709 15895
rect 26709 15861 26743 15895
rect 26743 15861 26752 15895
rect 26700 15852 26752 15861
rect 4182 15750 4234 15802
rect 4246 15750 4298 15802
rect 4310 15750 4362 15802
rect 4374 15750 4426 15802
rect 4438 15750 4490 15802
rect 4502 15750 4554 15802
rect 10182 15750 10234 15802
rect 10246 15750 10298 15802
rect 10310 15750 10362 15802
rect 10374 15750 10426 15802
rect 10438 15750 10490 15802
rect 10502 15750 10554 15802
rect 16182 15750 16234 15802
rect 16246 15750 16298 15802
rect 16310 15750 16362 15802
rect 16374 15750 16426 15802
rect 16438 15750 16490 15802
rect 16502 15750 16554 15802
rect 22182 15750 22234 15802
rect 22246 15750 22298 15802
rect 22310 15750 22362 15802
rect 22374 15750 22426 15802
rect 22438 15750 22490 15802
rect 22502 15750 22554 15802
rect 28182 15750 28234 15802
rect 28246 15750 28298 15802
rect 28310 15750 28362 15802
rect 28374 15750 28426 15802
rect 28438 15750 28490 15802
rect 28502 15750 28554 15802
rect 1860 15648 1912 15700
rect 4804 15648 4856 15700
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 6368 15648 6420 15700
rect 7840 15648 7892 15700
rect 10968 15648 11020 15700
rect 13176 15648 13228 15700
rect 13268 15648 13320 15700
rect 7932 15512 7984 15564
rect 2044 15444 2096 15453
rect 11612 15580 11664 15632
rect 10784 15512 10836 15564
rect 10876 15512 10928 15564
rect 15108 15648 15160 15700
rect 15384 15580 15436 15632
rect 16120 15580 16172 15632
rect 18328 15648 18380 15700
rect 19156 15648 19208 15700
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 4804 15376 4856 15428
rect 11428 15444 11480 15496
rect 5816 15376 5868 15428
rect 9588 15376 9640 15428
rect 7748 15308 7800 15360
rect 11888 15376 11940 15428
rect 12164 15444 12216 15496
rect 15568 15444 15620 15496
rect 18328 15444 18380 15496
rect 20904 15512 20956 15564
rect 22652 15648 22704 15700
rect 23848 15648 23900 15700
rect 26700 15648 26752 15700
rect 27528 15648 27580 15700
rect 25872 15512 25924 15564
rect 29644 15512 29696 15564
rect 17868 15376 17920 15428
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 10968 15308 11020 15360
rect 14096 15351 14148 15360
rect 14096 15317 14105 15351
rect 14105 15317 14139 15351
rect 14139 15317 14148 15351
rect 14096 15308 14148 15317
rect 15292 15351 15344 15360
rect 15292 15317 15301 15351
rect 15301 15317 15335 15351
rect 15335 15317 15344 15351
rect 15292 15308 15344 15317
rect 16212 15308 16264 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 18512 15376 18564 15428
rect 19248 15419 19300 15428
rect 19248 15385 19257 15419
rect 19257 15385 19291 15419
rect 19291 15385 19300 15419
rect 19248 15376 19300 15385
rect 19708 15444 19760 15496
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 26056 15487 26108 15496
rect 26056 15453 26065 15487
rect 26065 15453 26099 15487
rect 26099 15453 26108 15487
rect 26056 15444 26108 15453
rect 26516 15444 26568 15496
rect 20536 15308 20588 15360
rect 22008 15376 22060 15428
rect 24124 15376 24176 15428
rect 26976 15376 27028 15428
rect 27436 15376 27488 15428
rect 26700 15351 26752 15360
rect 26700 15317 26709 15351
rect 26709 15317 26743 15351
rect 26743 15317 26752 15351
rect 26700 15308 26752 15317
rect 27804 15351 27856 15360
rect 27804 15317 27813 15351
rect 27813 15317 27847 15351
rect 27847 15317 27856 15351
rect 27804 15308 27856 15317
rect 4922 15206 4974 15258
rect 4986 15206 5038 15258
rect 5050 15206 5102 15258
rect 5114 15206 5166 15258
rect 5178 15206 5230 15258
rect 5242 15206 5294 15258
rect 10922 15206 10974 15258
rect 10986 15206 11038 15258
rect 11050 15206 11102 15258
rect 11114 15206 11166 15258
rect 11178 15206 11230 15258
rect 11242 15206 11294 15258
rect 16922 15206 16974 15258
rect 16986 15206 17038 15258
rect 17050 15206 17102 15258
rect 17114 15206 17166 15258
rect 17178 15206 17230 15258
rect 17242 15206 17294 15258
rect 22922 15206 22974 15258
rect 22986 15206 23038 15258
rect 23050 15206 23102 15258
rect 23114 15206 23166 15258
rect 23178 15206 23230 15258
rect 23242 15206 23294 15258
rect 28922 15206 28974 15258
rect 28986 15206 29038 15258
rect 29050 15206 29102 15258
rect 29114 15206 29166 15258
rect 29178 15206 29230 15258
rect 29242 15206 29294 15258
rect 5816 15147 5868 15156
rect 5816 15113 5825 15147
rect 5825 15113 5859 15147
rect 5859 15113 5868 15147
rect 5816 15104 5868 15113
rect 6644 15104 6696 15156
rect 7840 15104 7892 15156
rect 7288 14968 7340 15020
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 9588 15147 9640 15156
rect 9588 15113 9597 15147
rect 9597 15113 9631 15147
rect 9631 15113 9640 15147
rect 9588 15104 9640 15113
rect 10692 15104 10744 15156
rect 12624 15104 12676 15156
rect 13176 15147 13228 15156
rect 13176 15113 13185 15147
rect 13185 15113 13219 15147
rect 13219 15113 13228 15147
rect 13176 15104 13228 15113
rect 14096 15104 14148 15156
rect 14464 15104 14516 15156
rect 15292 15104 15344 15156
rect 15936 15104 15988 15156
rect 18052 15104 18104 15156
rect 22008 15104 22060 15156
rect 26148 15104 26200 15156
rect 26700 15104 26752 15156
rect 8208 15079 8260 15088
rect 8208 15045 8217 15079
rect 8217 15045 8251 15079
rect 8251 15045 8260 15079
rect 8208 15036 8260 15045
rect 8484 14968 8536 15020
rect 11704 14968 11756 15020
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 6736 14832 6788 14884
rect 7288 14832 7340 14884
rect 8208 14832 8260 14884
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 13636 14900 13688 14952
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 12164 14764 12216 14816
rect 13728 14764 13780 14816
rect 15200 14968 15252 15020
rect 15568 15011 15620 15020
rect 15568 14977 15575 15011
rect 15575 14977 15620 15011
rect 15568 14968 15620 14977
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 16212 15036 16264 15088
rect 16120 15011 16172 15020
rect 16120 14977 16129 15011
rect 16129 14977 16163 15011
rect 16163 14977 16172 15011
rect 16120 14968 16172 14977
rect 14740 14900 14792 14952
rect 15292 14832 15344 14884
rect 17868 14900 17920 14952
rect 18512 14900 18564 14952
rect 20536 15011 20588 15020
rect 20536 14977 20545 15011
rect 20545 14977 20579 15011
rect 20579 14977 20588 15011
rect 20536 14968 20588 14977
rect 21916 14968 21968 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 22836 14968 22888 15020
rect 23848 14968 23900 15020
rect 25688 15011 25740 15020
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 26148 14968 26200 15020
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 27252 15104 27304 15156
rect 29644 15104 29696 15156
rect 26424 14968 26476 14977
rect 24308 14900 24360 14952
rect 26056 14900 26108 14952
rect 26332 14900 26384 14952
rect 27804 15036 27856 15088
rect 27160 14900 27212 14952
rect 17960 14832 18012 14884
rect 22008 14832 22060 14884
rect 26516 14832 26568 14884
rect 29368 14900 29420 14952
rect 17500 14807 17552 14816
rect 17500 14773 17509 14807
rect 17509 14773 17543 14807
rect 17543 14773 17552 14807
rect 17500 14764 17552 14773
rect 18972 14764 19024 14816
rect 19340 14764 19392 14816
rect 20628 14807 20680 14816
rect 20628 14773 20637 14807
rect 20637 14773 20671 14807
rect 20671 14773 20680 14807
rect 20628 14764 20680 14773
rect 24676 14764 24728 14816
rect 25872 14807 25924 14816
rect 25872 14773 25881 14807
rect 25881 14773 25915 14807
rect 25915 14773 25924 14807
rect 25872 14764 25924 14773
rect 26792 14764 26844 14816
rect 27252 14764 27304 14816
rect 4182 14662 4234 14714
rect 4246 14662 4298 14714
rect 4310 14662 4362 14714
rect 4374 14662 4426 14714
rect 4438 14662 4490 14714
rect 4502 14662 4554 14714
rect 10182 14662 10234 14714
rect 10246 14662 10298 14714
rect 10310 14662 10362 14714
rect 10374 14662 10426 14714
rect 10438 14662 10490 14714
rect 10502 14662 10554 14714
rect 16182 14662 16234 14714
rect 16246 14662 16298 14714
rect 16310 14662 16362 14714
rect 16374 14662 16426 14714
rect 16438 14662 16490 14714
rect 16502 14662 16554 14714
rect 22182 14662 22234 14714
rect 22246 14662 22298 14714
rect 22310 14662 22362 14714
rect 22374 14662 22426 14714
rect 22438 14662 22490 14714
rect 22502 14662 22554 14714
rect 28182 14662 28234 14714
rect 28246 14662 28298 14714
rect 28310 14662 28362 14714
rect 28374 14662 28426 14714
rect 28438 14662 28490 14714
rect 28502 14662 28554 14714
rect 11428 14560 11480 14612
rect 15292 14560 15344 14612
rect 15568 14603 15620 14612
rect 15568 14569 15577 14603
rect 15577 14569 15611 14603
rect 15611 14569 15620 14603
rect 15568 14560 15620 14569
rect 13912 14535 13964 14544
rect 13912 14501 13921 14535
rect 13921 14501 13955 14535
rect 13955 14501 13964 14535
rect 13912 14492 13964 14501
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 11888 14467 11940 14476
rect 11888 14433 11897 14467
rect 11897 14433 11931 14467
rect 11931 14433 11940 14467
rect 11888 14424 11940 14433
rect 13452 14424 13504 14476
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 17592 14560 17644 14612
rect 18512 14560 18564 14612
rect 26056 14560 26108 14612
rect 17500 14424 17552 14476
rect 26332 14424 26384 14476
rect 16856 14399 16908 14408
rect 16856 14365 16865 14399
rect 16865 14365 16899 14399
rect 16899 14365 16908 14399
rect 16856 14356 16908 14365
rect 26240 14356 26292 14408
rect 27160 14356 27212 14408
rect 13268 14220 13320 14272
rect 13636 14220 13688 14272
rect 13912 14288 13964 14340
rect 17868 14288 17920 14340
rect 27252 14288 27304 14340
rect 17960 14220 18012 14272
rect 4922 14118 4974 14170
rect 4986 14118 5038 14170
rect 5050 14118 5102 14170
rect 5114 14118 5166 14170
rect 5178 14118 5230 14170
rect 5242 14118 5294 14170
rect 10922 14118 10974 14170
rect 10986 14118 11038 14170
rect 11050 14118 11102 14170
rect 11114 14118 11166 14170
rect 11178 14118 11230 14170
rect 11242 14118 11294 14170
rect 16922 14118 16974 14170
rect 16986 14118 17038 14170
rect 17050 14118 17102 14170
rect 17114 14118 17166 14170
rect 17178 14118 17230 14170
rect 17242 14118 17294 14170
rect 22922 14118 22974 14170
rect 22986 14118 23038 14170
rect 23050 14118 23102 14170
rect 23114 14118 23166 14170
rect 23178 14118 23230 14170
rect 23242 14118 23294 14170
rect 28922 14118 28974 14170
rect 28986 14118 29038 14170
rect 29050 14118 29102 14170
rect 29114 14118 29166 14170
rect 29178 14118 29230 14170
rect 29242 14118 29294 14170
rect 3056 14059 3108 14068
rect 3056 14025 3065 14059
rect 3065 14025 3099 14059
rect 3099 14025 3108 14059
rect 3056 14016 3108 14025
rect 4068 14016 4120 14068
rect 8944 14016 8996 14068
rect 12440 14016 12492 14068
rect 12164 13991 12216 14000
rect 12164 13957 12173 13991
rect 12173 13957 12207 13991
rect 12207 13957 12216 13991
rect 12164 13948 12216 13957
rect 12256 13991 12308 14000
rect 12256 13957 12265 13991
rect 12265 13957 12299 13991
rect 12299 13957 12308 13991
rect 12256 13948 12308 13957
rect 12348 13948 12400 14000
rect 15752 14059 15804 14068
rect 15752 14025 15761 14059
rect 15761 14025 15795 14059
rect 15795 14025 15804 14059
rect 15752 14016 15804 14025
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 25504 14016 25556 14068
rect 2872 13880 2924 13932
rect 3240 13812 3292 13864
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 7840 13744 7892 13796
rect 8484 13744 8536 13796
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 12808 13880 12860 13932
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 18696 13948 18748 14000
rect 15108 13880 15160 13932
rect 14188 13812 14240 13864
rect 15752 13880 15804 13932
rect 24124 13880 24176 13932
rect 24400 13923 24452 13932
rect 24400 13889 24409 13923
rect 24409 13889 24443 13923
rect 24443 13889 24452 13923
rect 24400 13880 24452 13889
rect 24216 13812 24268 13864
rect 2228 13676 2280 13728
rect 2596 13719 2648 13728
rect 2596 13685 2605 13719
rect 2605 13685 2639 13719
rect 2639 13685 2648 13719
rect 2596 13676 2648 13685
rect 4160 13676 4212 13728
rect 8668 13676 8720 13728
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 21364 13676 21416 13728
rect 4182 13574 4234 13626
rect 4246 13574 4298 13626
rect 4310 13574 4362 13626
rect 4374 13574 4426 13626
rect 4438 13574 4490 13626
rect 4502 13574 4554 13626
rect 10182 13574 10234 13626
rect 10246 13574 10298 13626
rect 10310 13574 10362 13626
rect 10374 13574 10426 13626
rect 10438 13574 10490 13626
rect 10502 13574 10554 13626
rect 16182 13574 16234 13626
rect 16246 13574 16298 13626
rect 16310 13574 16362 13626
rect 16374 13574 16426 13626
rect 16438 13574 16490 13626
rect 16502 13574 16554 13626
rect 22182 13574 22234 13626
rect 22246 13574 22298 13626
rect 22310 13574 22362 13626
rect 22374 13574 22426 13626
rect 22438 13574 22490 13626
rect 22502 13574 22554 13626
rect 28182 13574 28234 13626
rect 28246 13574 28298 13626
rect 28310 13574 28362 13626
rect 28374 13574 28426 13626
rect 28438 13574 28490 13626
rect 28502 13574 28554 13626
rect 2596 13472 2648 13524
rect 2872 13472 2924 13524
rect 3976 13472 4028 13524
rect 4160 13472 4212 13524
rect 4528 13472 4580 13524
rect 4712 13472 4764 13524
rect 4620 13336 4672 13388
rect 2044 13268 2096 13320
rect 3792 13268 3844 13320
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6000 13311 6052 13320
rect 6000 13277 6007 13311
rect 6007 13277 6052 13311
rect 4712 13200 4764 13252
rect 6000 13268 6052 13277
rect 7748 13472 7800 13524
rect 9680 13472 9732 13524
rect 14096 13472 14148 13524
rect 15476 13472 15528 13524
rect 16120 13472 16172 13524
rect 9588 13404 9640 13456
rect 8668 13336 8720 13388
rect 9956 13336 10008 13388
rect 7288 13268 7340 13320
rect 7380 13311 7432 13320
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 9128 13268 9180 13320
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 6184 13243 6236 13252
rect 6184 13209 6193 13243
rect 6193 13209 6227 13243
rect 6227 13209 6236 13243
rect 6184 13200 6236 13209
rect 8208 13200 8260 13252
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 12900 13336 12952 13388
rect 20628 13404 20680 13456
rect 15844 13336 15896 13388
rect 25872 13472 25924 13524
rect 29368 13472 29420 13524
rect 11336 13268 11388 13320
rect 11888 13268 11940 13320
rect 14464 13268 14516 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 11520 13200 11572 13252
rect 14648 13200 14700 13252
rect 16120 13268 16172 13320
rect 22100 13268 22152 13320
rect 24676 13336 24728 13388
rect 23388 13268 23440 13320
rect 25780 13311 25832 13320
rect 25780 13277 25789 13311
rect 25789 13277 25823 13311
rect 25823 13277 25832 13311
rect 25780 13268 25832 13277
rect 18328 13200 18380 13252
rect 18604 13200 18656 13252
rect 19432 13200 19484 13252
rect 22376 13200 22428 13252
rect 22744 13200 22796 13252
rect 6460 13175 6512 13184
rect 6460 13141 6469 13175
rect 6469 13141 6503 13175
rect 6503 13141 6512 13175
rect 6460 13132 6512 13141
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 11336 13132 11388 13184
rect 15200 13132 15252 13184
rect 15844 13132 15896 13184
rect 21456 13132 21508 13184
rect 31300 13200 31352 13252
rect 24400 13175 24452 13184
rect 24400 13141 24409 13175
rect 24409 13141 24443 13175
rect 24443 13141 24452 13175
rect 24400 13132 24452 13141
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 4922 13030 4974 13082
rect 4986 13030 5038 13082
rect 5050 13030 5102 13082
rect 5114 13030 5166 13082
rect 5178 13030 5230 13082
rect 5242 13030 5294 13082
rect 10922 13030 10974 13082
rect 10986 13030 11038 13082
rect 11050 13030 11102 13082
rect 11114 13030 11166 13082
rect 11178 13030 11230 13082
rect 11242 13030 11294 13082
rect 16922 13030 16974 13082
rect 16986 13030 17038 13082
rect 17050 13030 17102 13082
rect 17114 13030 17166 13082
rect 17178 13030 17230 13082
rect 17242 13030 17294 13082
rect 22922 13030 22974 13082
rect 22986 13030 23038 13082
rect 23050 13030 23102 13082
rect 23114 13030 23166 13082
rect 23178 13030 23230 13082
rect 23242 13030 23294 13082
rect 28922 13030 28974 13082
rect 28986 13030 29038 13082
rect 29050 13030 29102 13082
rect 29114 13030 29166 13082
rect 29178 13030 29230 13082
rect 29242 13030 29294 13082
rect 2044 12792 2096 12844
rect 2228 12835 2280 12844
rect 2228 12801 2262 12835
rect 2262 12801 2280 12835
rect 2228 12792 2280 12801
rect 3792 12928 3844 12980
rect 3976 12928 4028 12980
rect 4712 12928 4764 12980
rect 5540 12928 5592 12980
rect 6000 12928 6052 12980
rect 5448 12860 5500 12912
rect 7196 12928 7248 12980
rect 7012 12860 7064 12912
rect 9036 12928 9088 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 9956 12928 10008 12980
rect 10692 12928 10744 12980
rect 10876 12928 10928 12980
rect 17316 12928 17368 12980
rect 18604 12928 18656 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 21088 12928 21140 12980
rect 21272 12928 21324 12980
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 7380 12860 7432 12912
rect 7932 12903 7984 12912
rect 7932 12869 7941 12903
rect 7941 12869 7975 12903
rect 7975 12869 7984 12903
rect 7932 12860 7984 12869
rect 4528 12724 4580 12776
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 5356 12792 5408 12844
rect 10508 12792 10560 12844
rect 6644 12724 6696 12776
rect 6828 12724 6880 12776
rect 10968 12860 11020 12912
rect 11612 12860 11664 12912
rect 14096 12860 14148 12912
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 19064 12835 19116 12844
rect 19064 12801 19073 12835
rect 19073 12801 19107 12835
rect 19107 12801 19116 12835
rect 19064 12792 19116 12801
rect 20352 12792 20404 12844
rect 23388 12928 23440 12980
rect 23480 12860 23532 12912
rect 24400 12928 24452 12980
rect 25228 12971 25280 12980
rect 25228 12937 25237 12971
rect 25237 12937 25271 12971
rect 25271 12937 25280 12971
rect 25228 12928 25280 12937
rect 25780 12928 25832 12980
rect 26424 12928 26476 12980
rect 29368 12928 29420 12980
rect 11152 12724 11204 12776
rect 11428 12724 11480 12776
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 17500 12724 17552 12776
rect 17776 12724 17828 12776
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 19800 12724 19852 12776
rect 20628 12767 20680 12776
rect 20628 12733 20637 12767
rect 20637 12733 20671 12767
rect 20671 12733 20680 12767
rect 21180 12835 21232 12844
rect 21180 12801 21194 12835
rect 21194 12801 21228 12835
rect 21228 12801 21232 12835
rect 21180 12792 21232 12801
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 21824 12835 21876 12844
rect 21824 12801 21833 12835
rect 21833 12801 21867 12835
rect 21867 12801 21876 12835
rect 21824 12792 21876 12801
rect 23204 12792 23256 12844
rect 24768 12860 24820 12912
rect 20628 12724 20680 12733
rect 6460 12656 6512 12708
rect 19708 12656 19760 12708
rect 23480 12724 23532 12776
rect 25872 12767 25924 12776
rect 25872 12733 25881 12767
rect 25881 12733 25915 12767
rect 25915 12733 25924 12767
rect 25872 12724 25924 12733
rect 26700 12767 26752 12776
rect 26700 12733 26709 12767
rect 26709 12733 26743 12767
rect 26743 12733 26752 12767
rect 26700 12724 26752 12733
rect 28080 12767 28132 12776
rect 28080 12733 28089 12767
rect 28089 12733 28123 12767
rect 28123 12733 28132 12767
rect 28080 12724 28132 12733
rect 5540 12588 5592 12640
rect 8852 12588 8904 12640
rect 11428 12588 11480 12640
rect 11704 12588 11756 12640
rect 11888 12588 11940 12640
rect 13728 12631 13780 12640
rect 13728 12597 13737 12631
rect 13737 12597 13771 12631
rect 13771 12597 13780 12631
rect 13728 12588 13780 12597
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 18696 12588 18748 12640
rect 20720 12588 20772 12640
rect 22744 12588 22796 12640
rect 23112 12588 23164 12640
rect 23664 12588 23716 12640
rect 26424 12588 26476 12640
rect 28632 12588 28684 12640
rect 4182 12486 4234 12538
rect 4246 12486 4298 12538
rect 4310 12486 4362 12538
rect 4374 12486 4426 12538
rect 4438 12486 4490 12538
rect 4502 12486 4554 12538
rect 10182 12486 10234 12538
rect 10246 12486 10298 12538
rect 10310 12486 10362 12538
rect 10374 12486 10426 12538
rect 10438 12486 10490 12538
rect 10502 12486 10554 12538
rect 16182 12486 16234 12538
rect 16246 12486 16298 12538
rect 16310 12486 16362 12538
rect 16374 12486 16426 12538
rect 16438 12486 16490 12538
rect 16502 12486 16554 12538
rect 22182 12486 22234 12538
rect 22246 12486 22298 12538
rect 22310 12486 22362 12538
rect 22374 12486 22426 12538
rect 22438 12486 22490 12538
rect 22502 12486 22554 12538
rect 28182 12486 28234 12538
rect 28246 12486 28298 12538
rect 28310 12486 28362 12538
rect 28374 12486 28426 12538
rect 28438 12486 28490 12538
rect 28502 12486 28554 12538
rect 5448 12384 5500 12436
rect 7932 12384 7984 12436
rect 8208 12427 8260 12436
rect 8208 12393 8217 12427
rect 8217 12393 8251 12427
rect 8251 12393 8260 12427
rect 8208 12384 8260 12393
rect 10600 12384 10652 12436
rect 10692 12384 10744 12436
rect 6184 12316 6236 12368
rect 6828 12248 6880 12300
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 8944 12316 8996 12368
rect 10508 12316 10560 12368
rect 11336 12384 11388 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 17040 12384 17092 12436
rect 8852 12180 8904 12232
rect 13452 12316 13504 12368
rect 5540 12112 5592 12164
rect 4712 12044 4764 12096
rect 5448 12044 5500 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 10692 12223 10744 12232
rect 10692 12189 10702 12223
rect 10702 12189 10736 12223
rect 10736 12189 10744 12223
rect 10692 12180 10744 12189
rect 10416 12112 10468 12164
rect 9680 12044 9732 12096
rect 10784 12044 10836 12096
rect 11060 12044 11112 12096
rect 12072 12180 12124 12232
rect 12256 12223 12308 12232
rect 12256 12189 12265 12223
rect 12265 12189 12299 12223
rect 12299 12189 12308 12223
rect 12256 12180 12308 12189
rect 13728 12248 13780 12300
rect 17408 12248 17460 12300
rect 17684 12248 17736 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 21732 12384 21784 12436
rect 23572 12384 23624 12436
rect 23664 12384 23716 12436
rect 24032 12384 24084 12436
rect 24216 12427 24268 12436
rect 24216 12393 24225 12427
rect 24225 12393 24259 12427
rect 24259 12393 24268 12427
rect 24216 12384 24268 12393
rect 23204 12316 23256 12368
rect 26700 12384 26752 12436
rect 30656 12384 30708 12436
rect 15384 12180 15436 12232
rect 17592 12180 17644 12232
rect 14188 12112 14240 12164
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 19340 12112 19392 12164
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 21732 12155 21784 12164
rect 21732 12121 21766 12155
rect 21766 12121 21784 12155
rect 11612 12044 11664 12096
rect 12072 12087 12124 12096
rect 12072 12053 12081 12087
rect 12081 12053 12115 12087
rect 12115 12053 12124 12087
rect 12072 12044 12124 12053
rect 12716 12044 12768 12096
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 17868 12044 17920 12096
rect 18052 12044 18104 12096
rect 19432 12044 19484 12096
rect 21732 12112 21784 12121
rect 23388 12180 23440 12232
rect 20996 12087 21048 12096
rect 20996 12053 21005 12087
rect 21005 12053 21039 12087
rect 21039 12053 21048 12087
rect 20996 12044 21048 12053
rect 23112 12155 23164 12164
rect 23112 12121 23121 12155
rect 23121 12121 23155 12155
rect 23155 12121 23164 12155
rect 23112 12112 23164 12121
rect 23388 12044 23440 12096
rect 26240 12248 26292 12300
rect 23572 12044 23624 12096
rect 24308 12180 24360 12232
rect 24492 12180 24544 12232
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 26608 12180 26660 12232
rect 26700 12223 26752 12232
rect 26700 12189 26709 12223
rect 26709 12189 26743 12223
rect 26743 12189 26752 12223
rect 26700 12180 26752 12189
rect 26976 12180 27028 12232
rect 24216 12112 24268 12164
rect 26148 12112 26200 12164
rect 27620 12155 27672 12164
rect 27620 12121 27629 12155
rect 27629 12121 27663 12155
rect 27663 12121 27672 12155
rect 27620 12112 27672 12121
rect 28632 12112 28684 12164
rect 25228 12044 25280 12096
rect 26884 12087 26936 12096
rect 26884 12053 26893 12087
rect 26893 12053 26927 12087
rect 26927 12053 26936 12087
rect 26884 12044 26936 12053
rect 4922 11942 4974 11994
rect 4986 11942 5038 11994
rect 5050 11942 5102 11994
rect 5114 11942 5166 11994
rect 5178 11942 5230 11994
rect 5242 11942 5294 11994
rect 10922 11942 10974 11994
rect 10986 11942 11038 11994
rect 11050 11942 11102 11994
rect 11114 11942 11166 11994
rect 11178 11942 11230 11994
rect 11242 11942 11294 11994
rect 16922 11942 16974 11994
rect 16986 11942 17038 11994
rect 17050 11942 17102 11994
rect 17114 11942 17166 11994
rect 17178 11942 17230 11994
rect 17242 11942 17294 11994
rect 22922 11942 22974 11994
rect 22986 11942 23038 11994
rect 23050 11942 23102 11994
rect 23114 11942 23166 11994
rect 23178 11942 23230 11994
rect 23242 11942 23294 11994
rect 28922 11942 28974 11994
rect 28986 11942 29038 11994
rect 29050 11942 29102 11994
rect 29114 11942 29166 11994
rect 29178 11942 29230 11994
rect 29242 11942 29294 11994
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 6552 11840 6604 11892
rect 940 11704 992 11756
rect 4804 11704 4856 11756
rect 10508 11840 10560 11892
rect 10876 11840 10928 11892
rect 12072 11840 12124 11892
rect 13820 11840 13872 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 14188 11840 14240 11849
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 9588 11704 9640 11756
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 9772 11704 9824 11756
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 9680 11568 9732 11620
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 14832 11704 14884 11756
rect 11888 11568 11940 11620
rect 12256 11568 12308 11620
rect 12900 11568 12952 11620
rect 14096 11568 14148 11620
rect 9956 11500 10008 11552
rect 10416 11500 10468 11552
rect 11796 11500 11848 11552
rect 12532 11500 12584 11552
rect 13176 11500 13228 11552
rect 16028 11704 16080 11756
rect 16672 11840 16724 11892
rect 18144 11840 18196 11892
rect 19064 11840 19116 11892
rect 21456 11840 21508 11892
rect 21732 11840 21784 11892
rect 15292 11636 15344 11688
rect 16580 11704 16632 11756
rect 16764 11772 16816 11824
rect 21916 11772 21968 11824
rect 23480 11840 23532 11892
rect 24492 11840 24544 11892
rect 14280 11568 14332 11620
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 17316 11500 17368 11552
rect 18052 11704 18104 11756
rect 18236 11704 18288 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18604 11704 18656 11756
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 20996 11704 21048 11756
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 21548 11704 21600 11756
rect 23388 11747 23440 11756
rect 23388 11713 23397 11747
rect 23397 11713 23431 11747
rect 23431 11713 23440 11747
rect 23388 11704 23440 11713
rect 26424 11840 26476 11892
rect 28080 11840 28132 11892
rect 26424 11747 26476 11756
rect 26424 11713 26433 11747
rect 26433 11713 26467 11747
rect 26467 11713 26476 11747
rect 26424 11704 26476 11713
rect 20444 11568 20496 11620
rect 30656 11704 30708 11756
rect 22652 11500 22704 11552
rect 26332 11500 26384 11552
rect 26516 11500 26568 11552
rect 26976 11679 27028 11688
rect 26976 11645 26985 11679
rect 26985 11645 27019 11679
rect 27019 11645 27028 11679
rect 26976 11636 27028 11645
rect 27712 11500 27764 11552
rect 4182 11398 4234 11450
rect 4246 11398 4298 11450
rect 4310 11398 4362 11450
rect 4374 11398 4426 11450
rect 4438 11398 4490 11450
rect 4502 11398 4554 11450
rect 10182 11398 10234 11450
rect 10246 11398 10298 11450
rect 10310 11398 10362 11450
rect 10374 11398 10426 11450
rect 10438 11398 10490 11450
rect 10502 11398 10554 11450
rect 16182 11398 16234 11450
rect 16246 11398 16298 11450
rect 16310 11398 16362 11450
rect 16374 11398 16426 11450
rect 16438 11398 16490 11450
rect 16502 11398 16554 11450
rect 22182 11398 22234 11450
rect 22246 11398 22298 11450
rect 22310 11398 22362 11450
rect 22374 11398 22426 11450
rect 22438 11398 22490 11450
rect 22502 11398 22554 11450
rect 28182 11398 28234 11450
rect 28246 11398 28298 11450
rect 28310 11398 28362 11450
rect 28374 11398 28426 11450
rect 28438 11398 28490 11450
rect 28502 11398 28554 11450
rect 4436 11296 4488 11348
rect 4620 11296 4672 11348
rect 10692 11296 10744 11348
rect 11336 11296 11388 11348
rect 9956 11228 10008 11280
rect 14740 11296 14792 11348
rect 17316 11339 17368 11348
rect 17316 11305 17325 11339
rect 17325 11305 17359 11339
rect 17359 11305 17368 11339
rect 17316 11296 17368 11305
rect 18328 11296 18380 11348
rect 18696 11296 18748 11348
rect 21456 11296 21508 11348
rect 26424 11296 26476 11348
rect 26792 11296 26844 11348
rect 26884 11296 26936 11348
rect 27620 11296 27672 11348
rect 27712 11296 27764 11348
rect 17868 11228 17920 11280
rect 2044 11160 2096 11212
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 7932 11160 7984 11212
rect 10876 11160 10928 11212
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 12532 11160 12584 11212
rect 20352 11160 20404 11212
rect 4712 11092 4764 11144
rect 8760 11092 8812 11144
rect 9588 11092 9640 11144
rect 2964 11024 3016 11076
rect 4620 11024 4672 11076
rect 11428 11024 11480 11076
rect 11796 11024 11848 11076
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 15108 11092 15160 11144
rect 16764 11092 16816 11144
rect 17224 11092 17276 11144
rect 12716 11024 12768 11076
rect 16028 11024 16080 11076
rect 19340 11024 19392 11076
rect 21548 11024 21600 11076
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 11612 10956 11664 11008
rect 12072 10956 12124 11008
rect 22652 11228 22704 11280
rect 22376 11092 22428 11144
rect 27160 11092 27212 11144
rect 27344 11092 27396 11144
rect 22376 10956 22428 11008
rect 25780 11024 25832 11076
rect 4922 10854 4974 10906
rect 4986 10854 5038 10906
rect 5050 10854 5102 10906
rect 5114 10854 5166 10906
rect 5178 10854 5230 10906
rect 5242 10854 5294 10906
rect 10922 10854 10974 10906
rect 10986 10854 11038 10906
rect 11050 10854 11102 10906
rect 11114 10854 11166 10906
rect 11178 10854 11230 10906
rect 11242 10854 11294 10906
rect 16922 10854 16974 10906
rect 16986 10854 17038 10906
rect 17050 10854 17102 10906
rect 17114 10854 17166 10906
rect 17178 10854 17230 10906
rect 17242 10854 17294 10906
rect 22922 10854 22974 10906
rect 22986 10854 23038 10906
rect 23050 10854 23102 10906
rect 23114 10854 23166 10906
rect 23178 10854 23230 10906
rect 23242 10854 23294 10906
rect 28922 10854 28974 10906
rect 28986 10854 29038 10906
rect 29050 10854 29102 10906
rect 29114 10854 29166 10906
rect 29178 10854 29230 10906
rect 29242 10854 29294 10906
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 4712 10795 4764 10804
rect 4712 10761 4721 10795
rect 4721 10761 4755 10795
rect 4755 10761 4764 10795
rect 4712 10752 4764 10761
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 5632 10752 5684 10804
rect 9680 10752 9732 10804
rect 25780 10752 25832 10804
rect 3792 10684 3844 10736
rect 4068 10684 4120 10736
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3976 10616 4028 10668
rect 3240 10548 3292 10600
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 10692 10616 10744 10668
rect 23848 10616 23900 10668
rect 6920 10548 6972 10600
rect 24492 10591 24544 10600
rect 24492 10557 24501 10591
rect 24501 10557 24535 10591
rect 24535 10557 24544 10591
rect 24492 10548 24544 10557
rect 4528 10480 4580 10532
rect 4804 10480 4856 10532
rect 4436 10412 4488 10464
rect 4896 10412 4948 10464
rect 21916 10412 21968 10464
rect 4182 10310 4234 10362
rect 4246 10310 4298 10362
rect 4310 10310 4362 10362
rect 4374 10310 4426 10362
rect 4438 10310 4490 10362
rect 4502 10310 4554 10362
rect 10182 10310 10234 10362
rect 10246 10310 10298 10362
rect 10310 10310 10362 10362
rect 10374 10310 10426 10362
rect 10438 10310 10490 10362
rect 10502 10310 10554 10362
rect 16182 10310 16234 10362
rect 16246 10310 16298 10362
rect 16310 10310 16362 10362
rect 16374 10310 16426 10362
rect 16438 10310 16490 10362
rect 16502 10310 16554 10362
rect 22182 10310 22234 10362
rect 22246 10310 22298 10362
rect 22310 10310 22362 10362
rect 22374 10310 22426 10362
rect 22438 10310 22490 10362
rect 22502 10310 22554 10362
rect 28182 10310 28234 10362
rect 28246 10310 28298 10362
rect 28310 10310 28362 10362
rect 28374 10310 28426 10362
rect 28438 10310 28490 10362
rect 28502 10310 28554 10362
rect 3148 10208 3200 10260
rect 4068 10208 4120 10260
rect 5448 10208 5500 10260
rect 23572 10208 23624 10260
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 4620 10004 4672 10056
rect 4712 10004 4764 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 4896 10004 4948 10056
rect 19432 10072 19484 10124
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 22560 10072 22612 10124
rect 5356 10004 5408 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9956 10004 10008 10056
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 22376 10004 22428 10056
rect 24952 10072 25004 10124
rect 25044 10004 25096 10056
rect 4804 9868 4856 9920
rect 22744 9936 22796 9988
rect 23572 9936 23624 9988
rect 6368 9868 6420 9920
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 19340 9868 19392 9920
rect 19616 9868 19668 9920
rect 23480 9911 23532 9920
rect 23480 9877 23489 9911
rect 23489 9877 23523 9911
rect 23523 9877 23532 9911
rect 23480 9868 23532 9877
rect 24216 9868 24268 9920
rect 24584 9868 24636 9920
rect 24860 9868 24912 9920
rect 25412 9911 25464 9920
rect 25412 9877 25421 9911
rect 25421 9877 25455 9911
rect 25455 9877 25464 9911
rect 25412 9868 25464 9877
rect 4922 9766 4974 9818
rect 4986 9766 5038 9818
rect 5050 9766 5102 9818
rect 5114 9766 5166 9818
rect 5178 9766 5230 9818
rect 5242 9766 5294 9818
rect 10922 9766 10974 9818
rect 10986 9766 11038 9818
rect 11050 9766 11102 9818
rect 11114 9766 11166 9818
rect 11178 9766 11230 9818
rect 11242 9766 11294 9818
rect 16922 9766 16974 9818
rect 16986 9766 17038 9818
rect 17050 9766 17102 9818
rect 17114 9766 17166 9818
rect 17178 9766 17230 9818
rect 17242 9766 17294 9818
rect 22922 9766 22974 9818
rect 22986 9766 23038 9818
rect 23050 9766 23102 9818
rect 23114 9766 23166 9818
rect 23178 9766 23230 9818
rect 23242 9766 23294 9818
rect 28922 9766 28974 9818
rect 28986 9766 29038 9818
rect 29050 9766 29102 9818
rect 29114 9766 29166 9818
rect 29178 9766 29230 9818
rect 29242 9766 29294 9818
rect 7196 9664 7248 9716
rect 9864 9664 9916 9716
rect 17408 9664 17460 9716
rect 7104 9596 7156 9648
rect 7288 9596 7340 9648
rect 8300 9596 8352 9648
rect 15384 9596 15436 9648
rect 18328 9596 18380 9648
rect 19248 9596 19300 9648
rect 21916 9664 21968 9716
rect 22376 9664 22428 9716
rect 23388 9664 23440 9716
rect 3792 9528 3844 9580
rect 5724 9528 5776 9580
rect 6368 9528 6420 9580
rect 7564 9571 7616 9580
rect 7564 9537 7571 9571
rect 7571 9537 7616 9571
rect 7564 9528 7616 9537
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 7840 9571 7892 9580
rect 7840 9537 7854 9571
rect 7854 9537 7888 9571
rect 7888 9537 7892 9571
rect 7840 9528 7892 9537
rect 8484 9528 8536 9580
rect 11060 9528 11112 9580
rect 12164 9528 12216 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 4344 9392 4396 9444
rect 6828 9460 6880 9512
rect 3792 9324 3844 9376
rect 4712 9324 4764 9376
rect 6000 9324 6052 9376
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 9864 9460 9916 9512
rect 10048 9460 10100 9512
rect 10968 9460 11020 9512
rect 12348 9503 12400 9512
rect 12348 9469 12357 9503
rect 12357 9469 12391 9503
rect 12391 9469 12400 9503
rect 12348 9460 12400 9469
rect 19156 9528 19208 9580
rect 19892 9528 19944 9580
rect 20812 9571 20864 9580
rect 20812 9537 20822 9571
rect 20822 9537 20856 9571
rect 20856 9537 20864 9571
rect 20812 9528 20864 9537
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 21180 9571 21232 9580
rect 21180 9537 21194 9571
rect 21194 9537 21228 9571
rect 21228 9537 21232 9571
rect 21180 9528 21232 9537
rect 9312 9367 9364 9376
rect 9312 9333 9321 9367
rect 9321 9333 9355 9367
rect 9355 9333 9364 9367
rect 9312 9324 9364 9333
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 17316 9503 17368 9512
rect 17316 9469 17325 9503
rect 17325 9469 17359 9503
rect 17359 9469 17368 9503
rect 17316 9460 17368 9469
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 16028 9324 16080 9376
rect 16580 9324 16632 9376
rect 18236 9392 18288 9444
rect 19064 9503 19116 9512
rect 19064 9469 19073 9503
rect 19073 9469 19107 9503
rect 19107 9469 19116 9503
rect 19064 9460 19116 9469
rect 19248 9503 19300 9512
rect 19248 9469 19257 9503
rect 19257 9469 19291 9503
rect 19291 9469 19300 9503
rect 19248 9460 19300 9469
rect 20904 9460 20956 9512
rect 23756 9664 23808 9716
rect 23664 9596 23716 9648
rect 24492 9664 24544 9716
rect 24860 9664 24912 9716
rect 25412 9664 25464 9716
rect 23388 9571 23440 9580
rect 23388 9537 23397 9571
rect 23397 9537 23431 9571
rect 23431 9537 23440 9571
rect 23388 9528 23440 9537
rect 23480 9528 23532 9580
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 22008 9367 22060 9376
rect 22008 9333 22017 9367
rect 22017 9333 22051 9367
rect 22051 9333 22060 9367
rect 22008 9324 22060 9333
rect 24032 9571 24084 9580
rect 24032 9537 24041 9571
rect 24041 9537 24075 9571
rect 24075 9537 24084 9571
rect 24032 9528 24084 9537
rect 24124 9392 24176 9444
rect 24768 9528 24820 9580
rect 24400 9460 24452 9512
rect 25412 9503 25464 9512
rect 25412 9469 25421 9503
rect 25421 9469 25455 9503
rect 25455 9469 25464 9503
rect 25412 9460 25464 9469
rect 25872 9460 25924 9512
rect 30748 9528 30800 9580
rect 26424 9460 26476 9512
rect 24308 9392 24360 9444
rect 24860 9392 24912 9444
rect 24952 9392 25004 9444
rect 25596 9324 25648 9376
rect 26056 9367 26108 9376
rect 26056 9333 26065 9367
rect 26065 9333 26099 9367
rect 26099 9333 26108 9367
rect 26056 9324 26108 9333
rect 4182 9222 4234 9274
rect 4246 9222 4298 9274
rect 4310 9222 4362 9274
rect 4374 9222 4426 9274
rect 4438 9222 4490 9274
rect 4502 9222 4554 9274
rect 10182 9222 10234 9274
rect 10246 9222 10298 9274
rect 10310 9222 10362 9274
rect 10374 9222 10426 9274
rect 10438 9222 10490 9274
rect 10502 9222 10554 9274
rect 16182 9222 16234 9274
rect 16246 9222 16298 9274
rect 16310 9222 16362 9274
rect 16374 9222 16426 9274
rect 16438 9222 16490 9274
rect 16502 9222 16554 9274
rect 22182 9222 22234 9274
rect 22246 9222 22298 9274
rect 22310 9222 22362 9274
rect 22374 9222 22426 9274
rect 22438 9222 22490 9274
rect 22502 9222 22554 9274
rect 28182 9222 28234 9274
rect 28246 9222 28298 9274
rect 28310 9222 28362 9274
rect 28374 9222 28426 9274
rect 28438 9222 28490 9274
rect 28502 9222 28554 9274
rect 4712 9052 4764 9104
rect 2780 8916 2832 8968
rect 3332 8916 3384 8968
rect 6184 9120 6236 9172
rect 6644 9120 6696 9172
rect 6000 9027 6052 9036
rect 6000 8993 6009 9027
rect 6009 8993 6043 9027
rect 6043 8993 6052 9027
rect 6000 8984 6052 8993
rect 7748 9120 7800 9172
rect 9312 9120 9364 9172
rect 10968 9052 11020 9104
rect 12348 9120 12400 9172
rect 19156 9120 19208 9172
rect 19248 9120 19300 9172
rect 19616 9120 19668 9172
rect 2320 8848 2372 8900
rect 6552 8916 6604 8968
rect 7104 8916 7156 8968
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 10508 8984 10560 9036
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 4068 8823 4120 8832
rect 4068 8789 4077 8823
rect 4077 8789 4111 8823
rect 4111 8789 4120 8823
rect 4068 8780 4120 8789
rect 4620 8780 4672 8832
rect 5632 8823 5684 8832
rect 5632 8789 5641 8823
rect 5641 8789 5675 8823
rect 5675 8789 5684 8823
rect 5632 8780 5684 8789
rect 8668 8848 8720 8900
rect 11060 8984 11112 9036
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8852 8780 8904 8832
rect 9956 8848 10008 8900
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11336 8959 11388 8968
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 11428 8780 11480 8832
rect 12532 8984 12584 9036
rect 12072 8959 12124 8968
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 12072 8925 12086 8959
rect 12086 8925 12120 8959
rect 12120 8925 12124 8959
rect 12072 8916 12124 8925
rect 13820 8984 13872 9036
rect 21088 9120 21140 9172
rect 23388 9120 23440 9172
rect 24124 9120 24176 9172
rect 25044 9120 25096 9172
rect 25596 9120 25648 9172
rect 13360 8848 13412 8900
rect 15936 8916 15988 8968
rect 17960 8959 18012 8968
rect 14832 8848 14884 8900
rect 17960 8925 17969 8959
rect 17969 8925 18003 8959
rect 18003 8925 18012 8959
rect 17960 8916 18012 8925
rect 18328 8916 18380 8968
rect 11704 8780 11756 8832
rect 11796 8780 11848 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 16028 8780 16080 8832
rect 16672 8848 16724 8900
rect 17500 8848 17552 8900
rect 18236 8848 18288 8900
rect 19156 8916 19208 8968
rect 18052 8780 18104 8832
rect 18788 8780 18840 8832
rect 20168 8848 20220 8900
rect 21824 8848 21876 8900
rect 23388 8916 23440 8968
rect 22192 8848 22244 8900
rect 24032 9052 24084 9104
rect 24584 9052 24636 9104
rect 24768 9052 24820 9104
rect 26056 9120 26108 9172
rect 22100 8780 22152 8832
rect 23480 8823 23532 8832
rect 23480 8789 23489 8823
rect 23489 8789 23523 8823
rect 23523 8789 23532 8823
rect 23480 8780 23532 8789
rect 24032 8823 24084 8832
rect 24032 8789 24041 8823
rect 24041 8789 24075 8823
rect 24075 8789 24084 8823
rect 24032 8780 24084 8789
rect 25780 8780 25832 8832
rect 25872 8780 25924 8832
rect 4922 8678 4974 8730
rect 4986 8678 5038 8730
rect 5050 8678 5102 8730
rect 5114 8678 5166 8730
rect 5178 8678 5230 8730
rect 5242 8678 5294 8730
rect 10922 8678 10974 8730
rect 10986 8678 11038 8730
rect 11050 8678 11102 8730
rect 11114 8678 11166 8730
rect 11178 8678 11230 8730
rect 11242 8678 11294 8730
rect 16922 8678 16974 8730
rect 16986 8678 17038 8730
rect 17050 8678 17102 8730
rect 17114 8678 17166 8730
rect 17178 8678 17230 8730
rect 17242 8678 17294 8730
rect 22922 8678 22974 8730
rect 22986 8678 23038 8730
rect 23050 8678 23102 8730
rect 23114 8678 23166 8730
rect 23178 8678 23230 8730
rect 23242 8678 23294 8730
rect 28922 8678 28974 8730
rect 28986 8678 29038 8730
rect 29050 8678 29102 8730
rect 29114 8678 29166 8730
rect 29178 8678 29230 8730
rect 29242 8678 29294 8730
rect 2780 8508 2832 8560
rect 4068 8576 4120 8628
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 7564 8576 7616 8628
rect 4620 8508 4672 8560
rect 2688 8483 2740 8492
rect 2688 8449 2722 8483
rect 2722 8449 2740 8483
rect 2688 8440 2740 8449
rect 3976 8372 4028 8424
rect 4068 8372 4120 8424
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 4804 8440 4856 8492
rect 5356 8440 5408 8492
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 7932 8576 7984 8628
rect 8668 8440 8720 8492
rect 8852 8483 8904 8492
rect 8852 8449 8886 8483
rect 8886 8449 8904 8483
rect 8852 8440 8904 8449
rect 9220 8576 9272 8628
rect 11520 8576 11572 8628
rect 11796 8576 11848 8628
rect 10508 8440 10560 8492
rect 12164 8576 12216 8628
rect 13360 8619 13412 8628
rect 13360 8585 13369 8619
rect 13369 8585 13403 8619
rect 13403 8585 13412 8619
rect 13360 8576 13412 8585
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 3792 8304 3844 8356
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 9956 8347 10008 8356
rect 9956 8313 9965 8347
rect 9965 8313 9999 8347
rect 9999 8313 10008 8347
rect 9956 8304 10008 8313
rect 12532 8440 12584 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 15476 8576 15528 8628
rect 13544 8372 13596 8424
rect 14372 8372 14424 8424
rect 16580 8440 16632 8492
rect 17960 8440 18012 8492
rect 19064 8576 19116 8628
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 19892 8576 19944 8628
rect 20168 8576 20220 8628
rect 21088 8576 21140 8628
rect 21824 8576 21876 8628
rect 22008 8576 22060 8628
rect 23480 8576 23532 8628
rect 24952 8576 25004 8628
rect 25780 8576 25832 8628
rect 18696 8551 18748 8560
rect 18696 8517 18705 8551
rect 18705 8517 18739 8551
rect 18739 8517 18748 8551
rect 18696 8508 18748 8517
rect 18788 8551 18840 8560
rect 18788 8517 18797 8551
rect 18797 8517 18831 8551
rect 18831 8517 18840 8551
rect 18788 8508 18840 8517
rect 18604 8440 18656 8492
rect 7012 8236 7064 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 16488 8372 16540 8424
rect 16672 8304 16724 8356
rect 19800 8372 19852 8424
rect 24032 8440 24084 8492
rect 25872 8440 25924 8492
rect 22100 8415 22152 8424
rect 22100 8381 22109 8415
rect 22109 8381 22143 8415
rect 22143 8381 22152 8415
rect 22100 8372 22152 8381
rect 23572 8372 23624 8424
rect 15016 8279 15068 8288
rect 15016 8245 15025 8279
rect 15025 8245 15059 8279
rect 15059 8245 15068 8279
rect 15016 8236 15068 8245
rect 4182 8134 4234 8186
rect 4246 8134 4298 8186
rect 4310 8134 4362 8186
rect 4374 8134 4426 8186
rect 4438 8134 4490 8186
rect 4502 8134 4554 8186
rect 10182 8134 10234 8186
rect 10246 8134 10298 8186
rect 10310 8134 10362 8186
rect 10374 8134 10426 8186
rect 10438 8134 10490 8186
rect 10502 8134 10554 8186
rect 16182 8134 16234 8186
rect 16246 8134 16298 8186
rect 16310 8134 16362 8186
rect 16374 8134 16426 8186
rect 16438 8134 16490 8186
rect 16502 8134 16554 8186
rect 22182 8134 22234 8186
rect 22246 8134 22298 8186
rect 22310 8134 22362 8186
rect 22374 8134 22426 8186
rect 22438 8134 22490 8186
rect 22502 8134 22554 8186
rect 28182 8134 28234 8186
rect 28246 8134 28298 8186
rect 28310 8134 28362 8186
rect 28374 8134 28426 8186
rect 28438 8134 28490 8186
rect 28502 8134 28554 8186
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 7104 8032 7156 8084
rect 12532 8032 12584 8084
rect 30748 8075 30800 8084
rect 30748 8041 30757 8075
rect 30757 8041 30791 8075
rect 30791 8041 30800 8075
rect 30748 8032 30800 8041
rect 15936 7964 15988 8016
rect 17316 7896 17368 7948
rect 3884 7828 3936 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 9864 7828 9916 7880
rect 11336 7828 11388 7880
rect 12164 7828 12216 7880
rect 14832 7828 14884 7880
rect 15016 7871 15068 7880
rect 15016 7837 15050 7871
rect 15050 7837 15068 7871
rect 15016 7828 15068 7837
rect 18328 8007 18380 8016
rect 18328 7973 18337 8007
rect 18337 7973 18371 8007
rect 18371 7973 18380 8007
rect 18328 7964 18380 7973
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 18604 7828 18656 7880
rect 18696 7828 18748 7880
rect 31300 7828 31352 7880
rect 16304 7692 16356 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 17868 7692 17920 7744
rect 21640 7692 21692 7744
rect 4922 7590 4974 7642
rect 4986 7590 5038 7642
rect 5050 7590 5102 7642
rect 5114 7590 5166 7642
rect 5178 7590 5230 7642
rect 5242 7590 5294 7642
rect 10922 7590 10974 7642
rect 10986 7590 11038 7642
rect 11050 7590 11102 7642
rect 11114 7590 11166 7642
rect 11178 7590 11230 7642
rect 11242 7590 11294 7642
rect 16922 7590 16974 7642
rect 16986 7590 17038 7642
rect 17050 7590 17102 7642
rect 17114 7590 17166 7642
rect 17178 7590 17230 7642
rect 17242 7590 17294 7642
rect 22922 7590 22974 7642
rect 22986 7590 23038 7642
rect 23050 7590 23102 7642
rect 23114 7590 23166 7642
rect 23178 7590 23230 7642
rect 23242 7590 23294 7642
rect 28922 7590 28974 7642
rect 28986 7590 29038 7642
rect 29050 7590 29102 7642
rect 29114 7590 29166 7642
rect 29178 7590 29230 7642
rect 29242 7590 29294 7642
rect 14648 7488 14700 7540
rect 16304 7531 16356 7540
rect 16304 7497 16313 7531
rect 16313 7497 16347 7531
rect 16347 7497 16356 7531
rect 16304 7488 16356 7497
rect 14832 7352 14884 7404
rect 4182 7046 4234 7098
rect 4246 7046 4298 7098
rect 4310 7046 4362 7098
rect 4374 7046 4426 7098
rect 4438 7046 4490 7098
rect 4502 7046 4554 7098
rect 10182 7046 10234 7098
rect 10246 7046 10298 7098
rect 10310 7046 10362 7098
rect 10374 7046 10426 7098
rect 10438 7046 10490 7098
rect 10502 7046 10554 7098
rect 16182 7046 16234 7098
rect 16246 7046 16298 7098
rect 16310 7046 16362 7098
rect 16374 7046 16426 7098
rect 16438 7046 16490 7098
rect 16502 7046 16554 7098
rect 22182 7046 22234 7098
rect 22246 7046 22298 7098
rect 22310 7046 22362 7098
rect 22374 7046 22426 7098
rect 22438 7046 22490 7098
rect 22502 7046 22554 7098
rect 28182 7046 28234 7098
rect 28246 7046 28298 7098
rect 28310 7046 28362 7098
rect 28374 7046 28426 7098
rect 28438 7046 28490 7098
rect 28502 7046 28554 7098
rect 5908 6740 5960 6792
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 6828 6808 6880 6860
rect 7932 6851 7984 6860
rect 7932 6817 7941 6851
rect 7941 6817 7975 6851
rect 7975 6817 7984 6851
rect 20996 6944 21048 6996
rect 7932 6808 7984 6817
rect 7012 6740 7064 6792
rect 8116 6783 8168 6792
rect 8116 6749 8126 6783
rect 8126 6749 8160 6783
rect 8160 6749 8168 6783
rect 8116 6740 8168 6749
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8484 6783 8536 6792
rect 8484 6749 8498 6783
rect 8498 6749 8532 6783
rect 8532 6749 8536 6783
rect 8484 6740 8536 6749
rect 11428 6740 11480 6792
rect 11520 6740 11572 6792
rect 18328 6740 18380 6792
rect 19800 6851 19852 6860
rect 19800 6817 19809 6851
rect 19809 6817 19843 6851
rect 19843 6817 19852 6851
rect 19800 6808 19852 6817
rect 10784 6672 10836 6724
rect 8024 6604 8076 6656
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 9680 6604 9732 6656
rect 9956 6647 10008 6656
rect 9956 6613 9965 6647
rect 9965 6613 9999 6647
rect 9999 6613 10008 6647
rect 9956 6604 10008 6613
rect 11336 6604 11388 6656
rect 19432 6740 19484 6792
rect 20720 6783 20772 6792
rect 19156 6604 19208 6656
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 19708 6647 19760 6656
rect 19708 6613 19717 6647
rect 19717 6613 19751 6647
rect 19751 6613 19760 6647
rect 19708 6604 19760 6613
rect 19800 6604 19852 6656
rect 20812 6604 20864 6656
rect 20996 6604 21048 6656
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 22652 6944 22704 6996
rect 22652 6740 22704 6792
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 22008 6604 22060 6656
rect 22468 6715 22520 6724
rect 22468 6681 22477 6715
rect 22477 6681 22511 6715
rect 22511 6681 22520 6715
rect 22468 6672 22520 6681
rect 22652 6604 22704 6656
rect 24308 6672 24360 6724
rect 24584 6740 24636 6792
rect 24860 6783 24912 6792
rect 24860 6749 24874 6783
rect 24874 6749 24908 6783
rect 24908 6749 24912 6783
rect 24860 6740 24912 6749
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 24768 6715 24820 6724
rect 24768 6681 24777 6715
rect 24777 6681 24811 6715
rect 24811 6681 24820 6715
rect 24768 6672 24820 6681
rect 26240 6604 26292 6656
rect 4922 6502 4974 6554
rect 4986 6502 5038 6554
rect 5050 6502 5102 6554
rect 5114 6502 5166 6554
rect 5178 6502 5230 6554
rect 5242 6502 5294 6554
rect 10922 6502 10974 6554
rect 10986 6502 11038 6554
rect 11050 6502 11102 6554
rect 11114 6502 11166 6554
rect 11178 6502 11230 6554
rect 11242 6502 11294 6554
rect 16922 6502 16974 6554
rect 16986 6502 17038 6554
rect 17050 6502 17102 6554
rect 17114 6502 17166 6554
rect 17178 6502 17230 6554
rect 17242 6502 17294 6554
rect 22922 6502 22974 6554
rect 22986 6502 23038 6554
rect 23050 6502 23102 6554
rect 23114 6502 23166 6554
rect 23178 6502 23230 6554
rect 23242 6502 23294 6554
rect 28922 6502 28974 6554
rect 28986 6502 29038 6554
rect 29050 6502 29102 6554
rect 29114 6502 29166 6554
rect 29178 6502 29230 6554
rect 29242 6502 29294 6554
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 6000 6400 6052 6452
rect 7932 6400 7984 6452
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 8668 6400 8720 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 9956 6400 10008 6452
rect 13820 6400 13872 6452
rect 19248 6400 19300 6452
rect 20720 6400 20772 6452
rect 21548 6400 21600 6452
rect 22468 6400 22520 6452
rect 23572 6400 23624 6452
rect 24216 6400 24268 6452
rect 24676 6400 24728 6452
rect 24768 6400 24820 6452
rect 4068 6128 4120 6180
rect 6184 6196 6236 6248
rect 6276 6196 6328 6248
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 6368 6128 6420 6180
rect 8944 6264 8996 6316
rect 10048 6264 10100 6316
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10600 6103 10652 6112
rect 10600 6069 10609 6103
rect 10609 6069 10643 6103
rect 10643 6069 10652 6103
rect 10600 6060 10652 6069
rect 11980 6264 12032 6316
rect 10784 6196 10836 6248
rect 11612 6239 11664 6248
rect 11612 6205 11621 6239
rect 11621 6205 11655 6239
rect 11655 6205 11664 6239
rect 11612 6196 11664 6205
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 18236 6307 18288 6316
rect 18236 6273 18270 6307
rect 18270 6273 18288 6307
rect 18236 6264 18288 6273
rect 22100 6332 22152 6384
rect 13820 6196 13872 6248
rect 15200 6239 15252 6248
rect 15200 6205 15209 6239
rect 15209 6205 15243 6239
rect 15243 6205 15252 6239
rect 15200 6196 15252 6205
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 24400 6264 24452 6316
rect 14188 6128 14240 6180
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 20444 6128 20496 6180
rect 19340 6103 19392 6112
rect 19340 6069 19349 6103
rect 19349 6069 19383 6103
rect 19383 6069 19392 6103
rect 22008 6196 22060 6248
rect 24308 6128 24360 6180
rect 25412 6128 25464 6180
rect 19340 6060 19392 6069
rect 22652 6103 22704 6112
rect 22652 6069 22661 6103
rect 22661 6069 22695 6103
rect 22695 6069 22704 6103
rect 22652 6060 22704 6069
rect 24124 6103 24176 6112
rect 24124 6069 24133 6103
rect 24133 6069 24167 6103
rect 24167 6069 24176 6103
rect 24124 6060 24176 6069
rect 24216 6103 24268 6112
rect 24216 6069 24225 6103
rect 24225 6069 24259 6103
rect 24259 6069 24268 6103
rect 24216 6060 24268 6069
rect 4182 5958 4234 6010
rect 4246 5958 4298 6010
rect 4310 5958 4362 6010
rect 4374 5958 4426 6010
rect 4438 5958 4490 6010
rect 4502 5958 4554 6010
rect 10182 5958 10234 6010
rect 10246 5958 10298 6010
rect 10310 5958 10362 6010
rect 10374 5958 10426 6010
rect 10438 5958 10490 6010
rect 10502 5958 10554 6010
rect 16182 5958 16234 6010
rect 16246 5958 16298 6010
rect 16310 5958 16362 6010
rect 16374 5958 16426 6010
rect 16438 5958 16490 6010
rect 16502 5958 16554 6010
rect 22182 5958 22234 6010
rect 22246 5958 22298 6010
rect 22310 5958 22362 6010
rect 22374 5958 22426 6010
rect 22438 5958 22490 6010
rect 22502 5958 22554 6010
rect 28182 5958 28234 6010
rect 28246 5958 28298 6010
rect 28310 5958 28362 6010
rect 28374 5958 28426 6010
rect 28438 5958 28490 6010
rect 28502 5958 28554 6010
rect 5356 5856 5408 5908
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6000 5856 6052 5908
rect 6368 5856 6420 5908
rect 8116 5856 8168 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9772 5856 9824 5908
rect 8024 5652 8076 5704
rect 10600 5856 10652 5908
rect 11612 5856 11664 5908
rect 13636 5856 13688 5908
rect 15200 5856 15252 5908
rect 18236 5856 18288 5908
rect 10692 5720 10744 5772
rect 13544 5720 13596 5772
rect 11336 5695 11388 5704
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 11428 5695 11480 5704
rect 11428 5661 11438 5695
rect 11438 5661 11472 5695
rect 11472 5661 11480 5695
rect 11428 5652 11480 5661
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 12072 5652 12124 5704
rect 10600 5584 10652 5636
rect 11704 5627 11756 5636
rect 11704 5593 11713 5627
rect 11713 5593 11747 5627
rect 11747 5593 11756 5627
rect 11704 5584 11756 5593
rect 20444 5788 20496 5840
rect 19984 5720 20036 5772
rect 14832 5652 14884 5704
rect 4068 5516 4120 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 10140 5516 10192 5568
rect 11520 5516 11572 5568
rect 20996 5695 21048 5704
rect 20996 5661 21030 5695
rect 21030 5661 21048 5695
rect 22008 5856 22060 5908
rect 23204 5856 23256 5908
rect 24124 5856 24176 5908
rect 24216 5856 24268 5908
rect 24768 5856 24820 5908
rect 20996 5652 21048 5661
rect 22100 5652 22152 5704
rect 25412 5788 25464 5840
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 22284 5584 22336 5636
rect 23388 5584 23440 5636
rect 25504 5652 25556 5704
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 22192 5516 22244 5568
rect 23572 5516 23624 5568
rect 23664 5559 23716 5568
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 24768 5584 24820 5636
rect 27068 5652 27120 5704
rect 4922 5414 4974 5466
rect 4986 5414 5038 5466
rect 5050 5414 5102 5466
rect 5114 5414 5166 5466
rect 5178 5414 5230 5466
rect 5242 5414 5294 5466
rect 10922 5414 10974 5466
rect 10986 5414 11038 5466
rect 11050 5414 11102 5466
rect 11114 5414 11166 5466
rect 11178 5414 11230 5466
rect 11242 5414 11294 5466
rect 16922 5414 16974 5466
rect 16986 5414 17038 5466
rect 17050 5414 17102 5466
rect 17114 5414 17166 5466
rect 17178 5414 17230 5466
rect 17242 5414 17294 5466
rect 22922 5414 22974 5466
rect 22986 5414 23038 5466
rect 23050 5414 23102 5466
rect 23114 5414 23166 5466
rect 23178 5414 23230 5466
rect 23242 5414 23294 5466
rect 28922 5414 28974 5466
rect 28986 5414 29038 5466
rect 29050 5414 29102 5466
rect 29114 5414 29166 5466
rect 29178 5414 29230 5466
rect 29242 5414 29294 5466
rect 10784 5312 10836 5364
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 12624 5312 12676 5364
rect 12072 5244 12124 5296
rect 12348 5244 12400 5296
rect 15292 5312 15344 5364
rect 8760 5176 8812 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 9312 5176 9364 5228
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 17776 5244 17828 5296
rect 11428 5108 11480 5160
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14372 5108 14424 5160
rect 15200 5176 15252 5228
rect 22192 5355 22244 5364
rect 22192 5321 22201 5355
rect 22201 5321 22235 5355
rect 22235 5321 22244 5355
rect 22192 5312 22244 5321
rect 22652 5312 22704 5364
rect 23388 5312 23440 5364
rect 24308 5355 24360 5364
rect 24308 5321 24317 5355
rect 24317 5321 24351 5355
rect 24351 5321 24360 5355
rect 24308 5312 24360 5321
rect 23664 5244 23716 5296
rect 25320 5176 25372 5228
rect 25504 5176 25556 5228
rect 26700 5176 26752 5228
rect 14924 5040 14976 5092
rect 22836 5108 22888 5160
rect 22284 5040 22336 5092
rect 27068 5108 27120 5160
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 13820 4972 13872 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14188 4972 14240 5024
rect 16580 4972 16632 5024
rect 17408 4972 17460 5024
rect 26608 4972 26660 5024
rect 27436 5015 27488 5024
rect 27436 4981 27445 5015
rect 27445 4981 27479 5015
rect 27479 4981 27488 5015
rect 27436 4972 27488 4981
rect 4182 4870 4234 4922
rect 4246 4870 4298 4922
rect 4310 4870 4362 4922
rect 4374 4870 4426 4922
rect 4438 4870 4490 4922
rect 4502 4870 4554 4922
rect 10182 4870 10234 4922
rect 10246 4870 10298 4922
rect 10310 4870 10362 4922
rect 10374 4870 10426 4922
rect 10438 4870 10490 4922
rect 10502 4870 10554 4922
rect 16182 4870 16234 4922
rect 16246 4870 16298 4922
rect 16310 4870 16362 4922
rect 16374 4870 16426 4922
rect 16438 4870 16490 4922
rect 16502 4870 16554 4922
rect 22182 4870 22234 4922
rect 22246 4870 22298 4922
rect 22310 4870 22362 4922
rect 22374 4870 22426 4922
rect 22438 4870 22490 4922
rect 22502 4870 22554 4922
rect 28182 4870 28234 4922
rect 28246 4870 28298 4922
rect 28310 4870 28362 4922
rect 28374 4870 28426 4922
rect 28438 4870 28490 4922
rect 28502 4870 28554 4922
rect 9312 4768 9364 4820
rect 9772 4700 9824 4752
rect 12624 4768 12676 4820
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 10048 4564 10100 4616
rect 10600 4564 10652 4616
rect 9680 4428 9732 4480
rect 10692 4428 10744 4480
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12532 4496 12584 4548
rect 14096 4768 14148 4820
rect 14924 4768 14976 4820
rect 13820 4700 13872 4752
rect 15936 4700 15988 4752
rect 16028 4632 16080 4684
rect 14188 4564 14240 4616
rect 14372 4564 14424 4616
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 12900 4428 12952 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 14924 4471 14976 4480
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 17776 4564 17828 4616
rect 27436 4768 27488 4820
rect 26240 4607 26292 4616
rect 26240 4573 26249 4607
rect 26249 4573 26283 4607
rect 26283 4573 26292 4607
rect 26240 4564 26292 4573
rect 27160 4564 27212 4616
rect 28724 4564 28776 4616
rect 18420 4496 18472 4548
rect 16672 4428 16724 4480
rect 17960 4428 18012 4480
rect 27620 4471 27672 4480
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 4922 4326 4974 4378
rect 4986 4326 5038 4378
rect 5050 4326 5102 4378
rect 5114 4326 5166 4378
rect 5178 4326 5230 4378
rect 5242 4326 5294 4378
rect 10922 4326 10974 4378
rect 10986 4326 11038 4378
rect 11050 4326 11102 4378
rect 11114 4326 11166 4378
rect 11178 4326 11230 4378
rect 11242 4326 11294 4378
rect 16922 4326 16974 4378
rect 16986 4326 17038 4378
rect 17050 4326 17102 4378
rect 17114 4326 17166 4378
rect 17178 4326 17230 4378
rect 17242 4326 17294 4378
rect 22922 4326 22974 4378
rect 22986 4326 23038 4378
rect 23050 4326 23102 4378
rect 23114 4326 23166 4378
rect 23178 4326 23230 4378
rect 23242 4326 23294 4378
rect 28922 4326 28974 4378
rect 28986 4326 29038 4378
rect 29050 4326 29102 4378
rect 29114 4326 29166 4378
rect 29178 4326 29230 4378
rect 29242 4326 29294 4378
rect 16672 4224 16724 4276
rect 18420 4267 18472 4276
rect 18420 4233 18429 4267
rect 18429 4233 18463 4267
rect 18463 4233 18472 4267
rect 18420 4224 18472 4233
rect 9220 4088 9272 4140
rect 9588 4131 9640 4140
rect 9588 4097 9622 4131
rect 9622 4097 9640 4131
rect 9588 4088 9640 4097
rect 14924 4156 14976 4208
rect 27712 4156 27764 4208
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12440 4088 12492 4140
rect 13820 4088 13872 4140
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 14832 4020 14884 4072
rect 11428 3952 11480 4004
rect 17132 4088 17184 4140
rect 17684 4088 17736 4140
rect 17960 4088 18012 4140
rect 25504 4088 25556 4140
rect 19432 4020 19484 4072
rect 27620 4020 27672 4072
rect 14372 3884 14424 3936
rect 15384 3884 15436 3936
rect 17684 3927 17736 3936
rect 17684 3893 17693 3927
rect 17693 3893 17727 3927
rect 17727 3893 17736 3927
rect 17684 3884 17736 3893
rect 28724 3927 28776 3936
rect 28724 3893 28733 3927
rect 28733 3893 28767 3927
rect 28767 3893 28776 3927
rect 28724 3884 28776 3893
rect 4182 3782 4234 3834
rect 4246 3782 4298 3834
rect 4310 3782 4362 3834
rect 4374 3782 4426 3834
rect 4438 3782 4490 3834
rect 4502 3782 4554 3834
rect 10182 3782 10234 3834
rect 10246 3782 10298 3834
rect 10310 3782 10362 3834
rect 10374 3782 10426 3834
rect 10438 3782 10490 3834
rect 10502 3782 10554 3834
rect 16182 3782 16234 3834
rect 16246 3782 16298 3834
rect 16310 3782 16362 3834
rect 16374 3782 16426 3834
rect 16438 3782 16490 3834
rect 16502 3782 16554 3834
rect 22182 3782 22234 3834
rect 22246 3782 22298 3834
rect 22310 3782 22362 3834
rect 22374 3782 22426 3834
rect 22438 3782 22490 3834
rect 22502 3782 22554 3834
rect 28182 3782 28234 3834
rect 28246 3782 28298 3834
rect 28310 3782 28362 3834
rect 28374 3782 28426 3834
rect 28438 3782 28490 3834
rect 28502 3782 28554 3834
rect 10692 3680 10744 3732
rect 11888 3680 11940 3732
rect 12532 3680 12584 3732
rect 9220 3544 9272 3596
rect 11704 3544 11756 3596
rect 12992 3544 13044 3596
rect 13912 3587 13964 3596
rect 13912 3553 13921 3587
rect 13921 3553 13955 3587
rect 13955 3553 13964 3587
rect 13912 3544 13964 3553
rect 14832 3544 14884 3596
rect 17132 3723 17184 3732
rect 17132 3689 17141 3723
rect 17141 3689 17175 3723
rect 17175 3689 17184 3723
rect 17132 3680 17184 3689
rect 27712 3680 27764 3732
rect 27344 3612 27396 3664
rect 17684 3544 17736 3596
rect 9772 3408 9824 3460
rect 15936 3408 15988 3460
rect 15384 3340 15436 3392
rect 19432 3340 19484 3392
rect 20260 3340 20312 3392
rect 4922 3238 4974 3290
rect 4986 3238 5038 3290
rect 5050 3238 5102 3290
rect 5114 3238 5166 3290
rect 5178 3238 5230 3290
rect 5242 3238 5294 3290
rect 10922 3238 10974 3290
rect 10986 3238 11038 3290
rect 11050 3238 11102 3290
rect 11114 3238 11166 3290
rect 11178 3238 11230 3290
rect 11242 3238 11294 3290
rect 16922 3238 16974 3290
rect 16986 3238 17038 3290
rect 17050 3238 17102 3290
rect 17114 3238 17166 3290
rect 17178 3238 17230 3290
rect 17242 3238 17294 3290
rect 22922 3238 22974 3290
rect 22986 3238 23038 3290
rect 23050 3238 23102 3290
rect 23114 3238 23166 3290
rect 23178 3238 23230 3290
rect 23242 3238 23294 3290
rect 28922 3238 28974 3290
rect 28986 3238 29038 3290
rect 29050 3238 29102 3290
rect 29114 3238 29166 3290
rect 29178 3238 29230 3290
rect 29242 3238 29294 3290
rect 4182 2694 4234 2746
rect 4246 2694 4298 2746
rect 4310 2694 4362 2746
rect 4374 2694 4426 2746
rect 4438 2694 4490 2746
rect 4502 2694 4554 2746
rect 10182 2694 10234 2746
rect 10246 2694 10298 2746
rect 10310 2694 10362 2746
rect 10374 2694 10426 2746
rect 10438 2694 10490 2746
rect 10502 2694 10554 2746
rect 16182 2694 16234 2746
rect 16246 2694 16298 2746
rect 16310 2694 16362 2746
rect 16374 2694 16426 2746
rect 16438 2694 16490 2746
rect 16502 2694 16554 2746
rect 22182 2694 22234 2746
rect 22246 2694 22298 2746
rect 22310 2694 22362 2746
rect 22374 2694 22426 2746
rect 22438 2694 22490 2746
rect 22502 2694 22554 2746
rect 28182 2694 28234 2746
rect 28246 2694 28298 2746
rect 28310 2694 28362 2746
rect 28374 2694 28426 2746
rect 28438 2694 28490 2746
rect 28502 2694 28554 2746
rect 9864 2592 9916 2644
rect 13360 2456 13412 2508
rect 13912 2388 13964 2440
rect 19156 2388 19208 2440
rect 20260 2388 20312 2440
rect 28724 2388 28776 2440
rect 20 2320 72 2372
rect 10876 2363 10928 2372
rect 10876 2329 10885 2363
rect 10885 2329 10919 2363
rect 10919 2329 10928 2363
rect 10876 2320 10928 2329
rect 13268 2320 13320 2372
rect 28540 2363 28592 2372
rect 28540 2329 28549 2363
rect 28549 2329 28583 2363
rect 28583 2329 28592 2363
rect 28540 2320 28592 2329
rect 5356 2295 5408 2304
rect 5356 2261 5365 2295
rect 5365 2261 5399 2295
rect 5399 2261 5408 2295
rect 5356 2252 5408 2261
rect 16764 2295 16816 2304
rect 16764 2261 16773 2295
rect 16773 2261 16807 2295
rect 16807 2261 16816 2295
rect 16764 2252 16816 2261
rect 22560 2252 22612 2304
rect 30840 2295 30892 2304
rect 30840 2261 30849 2295
rect 30849 2261 30883 2295
rect 30883 2261 30892 2295
rect 30840 2252 30892 2261
rect 4922 2150 4974 2202
rect 4986 2150 5038 2202
rect 5050 2150 5102 2202
rect 5114 2150 5166 2202
rect 5178 2150 5230 2202
rect 5242 2150 5294 2202
rect 10922 2150 10974 2202
rect 10986 2150 11038 2202
rect 11050 2150 11102 2202
rect 11114 2150 11166 2202
rect 11178 2150 11230 2202
rect 11242 2150 11294 2202
rect 16922 2150 16974 2202
rect 16986 2150 17038 2202
rect 17050 2150 17102 2202
rect 17114 2150 17166 2202
rect 17178 2150 17230 2202
rect 17242 2150 17294 2202
rect 22922 2150 22974 2202
rect 22986 2150 23038 2202
rect 23050 2150 23102 2202
rect 23114 2150 23166 2202
rect 23178 2150 23230 2202
rect 23242 2150 23294 2202
rect 28922 2150 28974 2202
rect 28986 2150 29038 2202
rect 29050 2150 29102 2202
rect 29114 2150 29166 2202
rect 29178 2150 29230 2202
rect 29242 2150 29294 2202
<< metal2 >>
rect 1306 33796 1362 34596
rect 7102 33796 7158 34596
rect 12254 33796 12310 34596
rect 18050 33796 18106 34596
rect 23846 33796 23902 34596
rect 29642 33796 29698 34596
rect 1320 31822 1348 33796
rect 4180 32124 4556 32133
rect 4236 32122 4260 32124
rect 4316 32122 4340 32124
rect 4396 32122 4420 32124
rect 4476 32122 4500 32124
rect 4236 32070 4246 32122
rect 4490 32070 4500 32122
rect 4236 32068 4260 32070
rect 4316 32068 4340 32070
rect 4396 32068 4420 32070
rect 4476 32068 4500 32070
rect 4180 32059 4556 32068
rect 7116 31822 7144 33796
rect 10180 32124 10556 32133
rect 10236 32122 10260 32124
rect 10316 32122 10340 32124
rect 10396 32122 10420 32124
rect 10476 32122 10500 32124
rect 10236 32070 10246 32122
rect 10490 32070 10500 32122
rect 10236 32068 10260 32070
rect 10316 32068 10340 32070
rect 10396 32068 10420 32070
rect 10476 32068 10500 32070
rect 10180 32059 10556 32068
rect 12268 31822 12296 33796
rect 16180 32124 16556 32133
rect 16236 32122 16260 32124
rect 16316 32122 16340 32124
rect 16396 32122 16420 32124
rect 16476 32122 16500 32124
rect 16236 32070 16246 32122
rect 16490 32070 16500 32122
rect 16236 32068 16260 32070
rect 16316 32068 16340 32070
rect 16396 32068 16420 32070
rect 16476 32068 16500 32070
rect 16180 32059 16556 32068
rect 18064 32026 18092 33796
rect 22180 32124 22556 32133
rect 22236 32122 22260 32124
rect 22316 32122 22340 32124
rect 22396 32122 22420 32124
rect 22476 32122 22500 32124
rect 22236 32070 22246 32122
rect 22490 32070 22500 32122
rect 22236 32068 22260 32070
rect 22316 32068 22340 32070
rect 22396 32068 22420 32070
rect 22476 32068 22500 32070
rect 22180 32059 22556 32068
rect 23860 32026 23888 33796
rect 28180 32124 28556 32133
rect 28236 32122 28260 32124
rect 28316 32122 28340 32124
rect 28396 32122 28420 32124
rect 28476 32122 28500 32124
rect 28236 32070 28246 32122
rect 28490 32070 28500 32122
rect 28236 32068 28260 32070
rect 28316 32068 28340 32070
rect 28396 32068 28420 32070
rect 28476 32068 28500 32070
rect 28180 32059 28556 32068
rect 18052 32020 18104 32026
rect 18052 31962 18104 31968
rect 23848 32020 23900 32026
rect 23848 31962 23900 31968
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 1308 31816 1360 31822
rect 1308 31758 1360 31764
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 18144 31816 18196 31822
rect 18144 31758 18196 31764
rect 940 30252 992 30258
rect 940 30194 992 30200
rect 952 30025 980 30194
rect 938 30016 994 30025
rect 938 29951 994 29960
rect 940 24132 992 24138
rect 940 24074 992 24080
rect 952 23905 980 24074
rect 938 23896 994 23905
rect 938 23831 994 23840
rect 1688 19718 1716 31758
rect 12532 31680 12584 31686
rect 12532 31622 12584 31628
rect 4920 31580 5296 31589
rect 4976 31578 5000 31580
rect 5056 31578 5080 31580
rect 5136 31578 5160 31580
rect 5216 31578 5240 31580
rect 4976 31526 4986 31578
rect 5230 31526 5240 31578
rect 4976 31524 5000 31526
rect 5056 31524 5080 31526
rect 5136 31524 5160 31526
rect 5216 31524 5240 31526
rect 4920 31515 5296 31524
rect 10920 31580 11296 31589
rect 10976 31578 11000 31580
rect 11056 31578 11080 31580
rect 11136 31578 11160 31580
rect 11216 31578 11240 31580
rect 10976 31526 10986 31578
rect 11230 31526 11240 31578
rect 10976 31524 11000 31526
rect 11056 31524 11080 31526
rect 11136 31524 11160 31526
rect 11216 31524 11240 31526
rect 10920 31515 11296 31524
rect 12544 31414 12572 31622
rect 16920 31580 17296 31589
rect 16976 31578 17000 31580
rect 17056 31578 17080 31580
rect 17136 31578 17160 31580
rect 17216 31578 17240 31580
rect 16976 31526 16986 31578
rect 17230 31526 17240 31578
rect 16976 31524 17000 31526
rect 17056 31524 17080 31526
rect 17136 31524 17160 31526
rect 17216 31524 17240 31526
rect 16920 31515 17296 31524
rect 12532 31408 12584 31414
rect 12532 31350 12584 31356
rect 8576 31272 8628 31278
rect 8576 31214 8628 31220
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 17960 31272 18012 31278
rect 17960 31214 18012 31220
rect 7012 31136 7064 31142
rect 7012 31078 7064 31084
rect 4180 31036 4556 31045
rect 4236 31034 4260 31036
rect 4316 31034 4340 31036
rect 4396 31034 4420 31036
rect 4476 31034 4500 31036
rect 4236 30982 4246 31034
rect 4490 30982 4500 31034
rect 4236 30980 4260 30982
rect 4316 30980 4340 30982
rect 4396 30980 4420 30982
rect 4476 30980 4500 30982
rect 4180 30971 4556 30980
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 4920 30492 5296 30501
rect 4976 30490 5000 30492
rect 5056 30490 5080 30492
rect 5136 30490 5160 30492
rect 5216 30490 5240 30492
rect 4976 30438 4986 30490
rect 5230 30438 5240 30490
rect 4976 30436 5000 30438
rect 5056 30436 5080 30438
rect 5136 30436 5160 30438
rect 5216 30436 5240 30438
rect 4920 30427 5296 30436
rect 5644 30394 5672 30670
rect 7024 30394 7052 31078
rect 7380 30728 7432 30734
rect 7380 30670 7432 30676
rect 5632 30388 5684 30394
rect 5632 30330 5684 30336
rect 7012 30388 7064 30394
rect 7012 30330 7064 30336
rect 6000 30116 6052 30122
rect 6000 30058 6052 30064
rect 4180 29948 4556 29957
rect 4236 29946 4260 29948
rect 4316 29946 4340 29948
rect 4396 29946 4420 29948
rect 4476 29946 4500 29948
rect 4236 29894 4246 29946
rect 4490 29894 4500 29946
rect 4236 29892 4260 29894
rect 4316 29892 4340 29894
rect 4396 29892 4420 29894
rect 4476 29892 4500 29894
rect 4180 29883 4556 29892
rect 4920 29404 5296 29413
rect 4976 29402 5000 29404
rect 5056 29402 5080 29404
rect 5136 29402 5160 29404
rect 5216 29402 5240 29404
rect 4976 29350 4986 29402
rect 5230 29350 5240 29402
rect 4976 29348 5000 29350
rect 5056 29348 5080 29350
rect 5136 29348 5160 29350
rect 5216 29348 5240 29350
rect 4920 29339 5296 29348
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 4180 28860 4556 28869
rect 4236 28858 4260 28860
rect 4316 28858 4340 28860
rect 4396 28858 4420 28860
rect 4476 28858 4500 28860
rect 4236 28806 4246 28858
rect 4490 28806 4500 28858
rect 4236 28804 4260 28806
rect 4316 28804 4340 28806
rect 4396 28804 4420 28806
rect 4476 28804 4500 28806
rect 4180 28795 4556 28804
rect 4920 28316 5296 28325
rect 4976 28314 5000 28316
rect 5056 28314 5080 28316
rect 5136 28314 5160 28316
rect 5216 28314 5240 28316
rect 4976 28262 4986 28314
rect 5230 28262 5240 28314
rect 4976 28260 5000 28262
rect 5056 28260 5080 28262
rect 5136 28260 5160 28262
rect 5216 28260 5240 28262
rect 4920 28251 5296 28260
rect 5552 28218 5580 28902
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 4620 28076 4672 28082
rect 4620 28018 4672 28024
rect 4180 27772 4556 27781
rect 4236 27770 4260 27772
rect 4316 27770 4340 27772
rect 4396 27770 4420 27772
rect 4476 27770 4500 27772
rect 4236 27718 4246 27770
rect 4490 27718 4500 27770
rect 4236 27716 4260 27718
rect 4316 27716 4340 27718
rect 4396 27716 4420 27718
rect 4476 27716 4500 27718
rect 4180 27707 4556 27716
rect 4632 27674 4660 28018
rect 6012 28014 6040 30058
rect 7392 29170 7420 30670
rect 8116 30660 8168 30666
rect 8116 30602 8168 30608
rect 8128 30394 8156 30602
rect 8588 30598 8616 31214
rect 9140 30598 9168 31214
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10180 31036 10556 31045
rect 10236 31034 10260 31036
rect 10316 31034 10340 31036
rect 10396 31034 10420 31036
rect 10476 31034 10500 31036
rect 10236 30982 10246 31034
rect 10490 30982 10500 31034
rect 10236 30980 10260 30982
rect 10316 30980 10340 30982
rect 10396 30980 10420 30982
rect 10476 30980 10500 30982
rect 10180 30971 10556 30980
rect 10416 30864 10468 30870
rect 10416 30806 10468 30812
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 9128 30592 9180 30598
rect 9128 30534 9180 30540
rect 8116 30388 8168 30394
rect 8116 30330 8168 30336
rect 8024 30252 8076 30258
rect 8024 30194 8076 30200
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 6092 29096 6144 29102
rect 6092 29038 6144 29044
rect 6000 28008 6052 28014
rect 6000 27950 6052 27956
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 5368 27470 5396 27814
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 4920 27228 5296 27237
rect 4976 27226 5000 27228
rect 5056 27226 5080 27228
rect 5136 27226 5160 27228
rect 5216 27226 5240 27228
rect 4976 27174 4986 27226
rect 5230 27174 5240 27226
rect 4976 27172 5000 27174
rect 5056 27172 5080 27174
rect 5136 27172 5160 27174
rect 5216 27172 5240 27174
rect 4920 27163 5296 27172
rect 4180 26684 4556 26693
rect 4236 26682 4260 26684
rect 4316 26682 4340 26684
rect 4396 26682 4420 26684
rect 4476 26682 4500 26684
rect 4236 26630 4246 26682
rect 4490 26630 4500 26682
rect 4236 26628 4260 26630
rect 4316 26628 4340 26630
rect 4396 26628 4420 26630
rect 4476 26628 4500 26630
rect 4180 26619 4556 26628
rect 4920 26140 5296 26149
rect 4976 26138 5000 26140
rect 5056 26138 5080 26140
rect 5136 26138 5160 26140
rect 5216 26138 5240 26140
rect 4976 26086 4986 26138
rect 5230 26086 5240 26138
rect 4976 26084 5000 26086
rect 5056 26084 5080 26086
rect 5136 26084 5160 26086
rect 5216 26084 5240 26086
rect 4920 26075 5296 26084
rect 5540 25832 5592 25838
rect 5540 25774 5592 25780
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4180 25596 4556 25605
rect 4236 25594 4260 25596
rect 4316 25594 4340 25596
rect 4396 25594 4420 25596
rect 4476 25594 4500 25596
rect 4236 25542 4246 25594
rect 4490 25542 4500 25594
rect 4236 25540 4260 25542
rect 4316 25540 4340 25542
rect 4396 25540 4420 25542
rect 4476 25540 4500 25542
rect 4180 25531 4556 25540
rect 4908 25498 4936 25638
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3988 24818 4016 25094
rect 4724 24954 4752 25230
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 4180 24508 4556 24517
rect 4236 24506 4260 24508
rect 4316 24506 4340 24508
rect 4396 24506 4420 24508
rect 4476 24506 4500 24508
rect 4236 24454 4246 24506
rect 4490 24454 4500 24506
rect 4236 24452 4260 24454
rect 4316 24452 4340 24454
rect 4396 24452 4420 24454
rect 4476 24452 4500 24454
rect 4180 24443 4556 24452
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1872 20330 1900 24074
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4180 23420 4556 23429
rect 4236 23418 4260 23420
rect 4316 23418 4340 23420
rect 4396 23418 4420 23420
rect 4476 23418 4500 23420
rect 4236 23366 4246 23418
rect 4490 23366 4500 23418
rect 4236 23364 4260 23366
rect 4316 23364 4340 23366
rect 4396 23364 4420 23366
rect 4476 23364 4500 23366
rect 4180 23355 4556 23364
rect 4632 23118 4660 23462
rect 4724 23322 4752 24890
rect 4816 24886 4844 25094
rect 4920 25052 5296 25061
rect 4976 25050 5000 25052
rect 5056 25050 5080 25052
rect 5136 25050 5160 25052
rect 5216 25050 5240 25052
rect 4976 24998 4986 25050
rect 5230 24998 5240 25050
rect 4976 24996 5000 24998
rect 5056 24996 5080 24998
rect 5136 24996 5160 24998
rect 5216 24996 5240 24998
rect 4920 24987 5296 24996
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4264 22778 4292 22918
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3896 20942 3924 22510
rect 4180 22332 4556 22341
rect 4236 22330 4260 22332
rect 4316 22330 4340 22332
rect 4396 22330 4420 22332
rect 4476 22330 4500 22332
rect 4236 22278 4246 22330
rect 4490 22278 4500 22330
rect 4236 22276 4260 22278
rect 4316 22276 4340 22278
rect 4396 22276 4420 22278
rect 4476 22276 4500 22278
rect 4180 22267 4556 22276
rect 4816 22094 4844 24822
rect 4920 23964 5296 23973
rect 4976 23962 5000 23964
rect 5056 23962 5080 23964
rect 5136 23962 5160 23964
rect 5216 23962 5240 23964
rect 4976 23910 4986 23962
rect 5230 23910 5240 23962
rect 4976 23908 5000 23910
rect 5056 23908 5080 23910
rect 5136 23908 5160 23910
rect 5216 23908 5240 23910
rect 4920 23899 5296 23908
rect 5368 23662 5396 25434
rect 5448 25220 5500 25226
rect 5448 25162 5500 25168
rect 5460 24954 5488 25162
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5552 24682 5580 25774
rect 6012 25498 6040 27950
rect 6104 27878 6132 29038
rect 6368 28960 6420 28966
rect 6368 28902 6420 28908
rect 6460 28960 6512 28966
rect 6460 28902 6512 28908
rect 6380 28490 6408 28902
rect 6368 28484 6420 28490
rect 6368 28426 6420 28432
rect 6472 28370 6500 28902
rect 7024 28762 7052 29106
rect 7012 28756 7064 28762
rect 7012 28698 7064 28704
rect 7392 28626 7420 29106
rect 7380 28620 7432 28626
rect 7380 28562 7432 28568
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 6380 28342 6500 28370
rect 6380 28218 6408 28342
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6552 28212 6604 28218
rect 6552 28154 6604 28160
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6104 27402 6132 27814
rect 6092 27396 6144 27402
rect 6092 27338 6144 27344
rect 6000 25492 6052 25498
rect 6000 25434 6052 25440
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 6104 24886 6132 25094
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6380 24698 6408 28154
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 6472 27674 6500 28018
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 6564 27334 6592 28154
rect 7392 28082 7420 28562
rect 7380 28076 7432 28082
rect 7380 28018 7432 28024
rect 7196 27668 7248 27674
rect 7196 27610 7248 27616
rect 7208 27470 7236 27610
rect 7196 27464 7248 27470
rect 7196 27406 7248 27412
rect 6552 27328 6604 27334
rect 6552 27270 6604 27276
rect 5540 24676 5592 24682
rect 6380 24670 6500 24698
rect 5540 24618 5592 24624
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5908 23656 5960 23662
rect 5908 23598 5960 23604
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5356 23044 5408 23050
rect 5356 22986 5408 22992
rect 4920 22876 5296 22885
rect 4976 22874 5000 22876
rect 5056 22874 5080 22876
rect 5136 22874 5160 22876
rect 5216 22874 5240 22876
rect 4976 22822 4986 22874
rect 5230 22822 5240 22874
rect 4976 22820 5000 22822
rect 5056 22820 5080 22822
rect 5136 22820 5160 22822
rect 5216 22820 5240 22822
rect 4920 22811 5296 22820
rect 5368 22778 5396 22986
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 4724 22066 4844 22094
rect 5724 22092 5776 22098
rect 4180 21244 4556 21253
rect 4236 21242 4260 21244
rect 4316 21242 4340 21244
rect 4396 21242 4420 21244
rect 4476 21242 4500 21244
rect 4236 21190 4246 21242
rect 4490 21190 4500 21242
rect 4236 21188 4260 21190
rect 4316 21188 4340 21190
rect 4396 21188 4420 21190
rect 4476 21188 4500 21190
rect 4180 21179 4556 21188
rect 3884 20936 3936 20942
rect 3884 20878 3936 20884
rect 4160 20868 4212 20874
rect 4160 20810 4212 20816
rect 4172 20602 4200 20810
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 4180 20156 4556 20165
rect 4236 20154 4260 20156
rect 4316 20154 4340 20156
rect 4396 20154 4420 20156
rect 4476 20154 4500 20156
rect 4236 20102 4246 20154
rect 4490 20102 4500 20154
rect 4236 20100 4260 20102
rect 4316 20100 4340 20102
rect 4396 20100 4420 20102
rect 4476 20100 4500 20102
rect 4180 20091 4556 20100
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2240 18426 2268 18702
rect 2608 18698 2636 19110
rect 3344 18970 3372 19314
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 3804 18426 3832 19110
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 1412 17921 1440 18226
rect 1398 17912 1454 17921
rect 2424 17882 2452 18226
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 1398 17847 1454 17856
rect 2412 17876 2464 17882
rect 2412 17818 2464 17824
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16182 2360 16390
rect 2320 16176 2372 16182
rect 2320 16118 2372 16124
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15706 1900 15846
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1964 15484 1992 15982
rect 2044 15496 2096 15502
rect 1964 15456 2044 15484
rect 2044 15438 2096 15444
rect 2056 13326 2084 15438
rect 3068 14074 3096 18022
rect 3252 16658 3280 18158
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3620 17678 3648 18022
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3896 16182 3924 16730
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3988 16046 4016 18770
rect 4080 18086 4108 19110
rect 4180 19068 4556 19077
rect 4236 19066 4260 19068
rect 4316 19066 4340 19068
rect 4396 19066 4420 19068
rect 4476 19066 4500 19068
rect 4236 19014 4246 19066
rect 4490 19014 4500 19066
rect 4236 19012 4260 19014
rect 4316 19012 4340 19014
rect 4396 19012 4420 19014
rect 4476 19012 4500 19014
rect 4180 19003 4556 19012
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18426 4292 18566
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4540 18358 4568 18906
rect 4632 18426 4660 19246
rect 4724 19174 4752 22066
rect 5724 22034 5776 22040
rect 4920 21788 5296 21797
rect 4976 21786 5000 21788
rect 5056 21786 5080 21788
rect 5136 21786 5160 21788
rect 5216 21786 5240 21788
rect 4976 21734 4986 21786
rect 5230 21734 5240 21786
rect 4976 21732 5000 21734
rect 5056 21732 5080 21734
rect 5136 21732 5160 21734
rect 5216 21732 5240 21734
rect 4920 21723 5296 21732
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5184 21146 5212 21286
rect 5460 21146 5488 21286
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 4816 20398 4844 20810
rect 5736 20806 5764 22034
rect 5920 21010 5948 23598
rect 6012 22506 6040 23598
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6196 22574 6224 22918
rect 6288 22778 6316 22918
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6380 22506 6408 22578
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 6368 22500 6420 22506
rect 6368 22442 6420 22448
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 4920 20700 5296 20709
rect 4976 20698 5000 20700
rect 5056 20698 5080 20700
rect 5136 20698 5160 20700
rect 5216 20698 5240 20700
rect 4976 20646 4986 20698
rect 5230 20646 5240 20698
rect 4976 20644 5000 20646
rect 5056 20644 5080 20646
rect 5136 20644 5160 20646
rect 5216 20644 5240 20646
rect 4920 20635 5296 20644
rect 5368 20602 5396 20742
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4724 18426 4752 18838
rect 4816 18766 4844 20334
rect 5552 20058 5580 20402
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 4920 19612 5296 19621
rect 4976 19610 5000 19612
rect 5056 19610 5080 19612
rect 5136 19610 5160 19612
rect 5216 19610 5240 19612
rect 4976 19558 4986 19610
rect 5230 19558 5240 19610
rect 4976 19556 5000 19558
rect 5056 19556 5080 19558
rect 5136 19556 5160 19558
rect 5216 19556 5240 19558
rect 4920 19547 5296 19556
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18834 5120 19246
rect 5080 18828 5132 18834
rect 5080 18770 5132 18776
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 4540 18170 4568 18294
rect 4540 18142 4752 18170
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4180 17980 4556 17989
rect 4236 17978 4260 17980
rect 4316 17978 4340 17980
rect 4396 17978 4420 17980
rect 4476 17978 4500 17980
rect 4236 17926 4246 17978
rect 4490 17926 4500 17978
rect 4236 17924 4260 17926
rect 4316 17924 4340 17926
rect 4396 17924 4420 17926
rect 4476 17924 4500 17926
rect 4180 17915 4556 17924
rect 4180 16892 4556 16901
rect 4236 16890 4260 16892
rect 4316 16890 4340 16892
rect 4396 16890 4420 16892
rect 4476 16890 4500 16892
rect 4236 16838 4246 16890
rect 4490 16838 4500 16890
rect 4236 16836 4260 16838
rect 4316 16836 4340 16838
rect 4396 16836 4420 16838
rect 4476 16836 4500 16838
rect 4180 16827 4556 16836
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16250 4384 16526
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12850 2084 13262
rect 2240 12850 2268 13670
rect 2608 13530 2636 13670
rect 2884 13530 2912 13874
rect 3252 13870 3280 15846
rect 4180 15804 4556 15813
rect 4236 15802 4260 15804
rect 4316 15802 4340 15804
rect 4396 15802 4420 15804
rect 4476 15802 4500 15804
rect 4236 15750 4246 15802
rect 4490 15750 4500 15802
rect 4236 15748 4260 15750
rect 4316 15748 4340 15750
rect 4396 15748 4420 15750
rect 4476 15748 4500 15750
rect 4180 15739 4556 15748
rect 4180 14716 4556 14725
rect 4236 14714 4260 14716
rect 4316 14714 4340 14716
rect 4396 14714 4420 14716
rect 4476 14714 4500 14716
rect 4236 14662 4246 14714
rect 4490 14662 4500 14714
rect 4236 14660 4260 14662
rect 4316 14660 4340 14662
rect 4396 14660 4420 14662
rect 4476 14660 4500 14662
rect 4180 14651 4556 14660
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 2056 11218 2084 12786
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2976 10810 3004 11018
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10266 3188 10610
rect 3252 10606 3280 13806
rect 3988 13530 4016 13806
rect 4080 13716 4108 14010
rect 4160 13728 4212 13734
rect 4080 13688 4160 13716
rect 3976 13524 4028 13530
rect 4080 13512 4108 13688
rect 4160 13670 4212 13676
rect 4180 13628 4556 13637
rect 4236 13626 4260 13628
rect 4316 13626 4340 13628
rect 4396 13626 4420 13628
rect 4476 13626 4500 13628
rect 4236 13574 4246 13626
rect 4490 13574 4500 13626
rect 4236 13572 4260 13574
rect 4316 13572 4340 13574
rect 4396 13572 4420 13574
rect 4476 13572 4500 13574
rect 4180 13563 4556 13572
rect 4160 13524 4212 13530
rect 4080 13484 4160 13512
rect 3976 13466 4028 13472
rect 4160 13466 4212 13472
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3804 12986 3832 13262
rect 3988 12986 4016 13466
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4540 12782 4568 13466
rect 4632 13394 4660 16594
rect 4724 16182 4752 18142
rect 4816 17746 4844 18702
rect 4920 18524 5296 18533
rect 4976 18522 5000 18524
rect 5056 18522 5080 18524
rect 5136 18522 5160 18524
rect 5216 18522 5240 18524
rect 4976 18470 4986 18522
rect 5230 18470 5240 18522
rect 4976 18468 5000 18470
rect 5056 18468 5080 18470
rect 5136 18468 5160 18470
rect 5216 18468 5240 18470
rect 4920 18459 5296 18468
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 17882 5488 18226
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4920 17436 5296 17445
rect 4976 17434 5000 17436
rect 5056 17434 5080 17436
rect 5136 17434 5160 17436
rect 5216 17434 5240 17436
rect 4976 17382 4986 17434
rect 5230 17382 5240 17434
rect 4976 17380 5000 17382
rect 5056 17380 5080 17382
rect 5136 17380 5160 17382
rect 5216 17380 5240 17382
rect 4920 17371 5296 17380
rect 4920 16348 5296 16357
rect 4976 16346 5000 16348
rect 5056 16346 5080 16348
rect 5136 16346 5160 16348
rect 5216 16346 5240 16348
rect 4976 16294 4986 16346
rect 5230 16294 5240 16346
rect 4976 16292 5000 16294
rect 5056 16292 5080 16294
rect 5136 16292 5160 16294
rect 5216 16292 5240 16294
rect 4920 16283 5296 16292
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4724 13530 4752 16118
rect 5460 16114 5488 17818
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15706 4844 15846
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12866 4660 13330
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4724 12986 4752 13194
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4632 12838 4752 12866
rect 4816 12850 4844 15370
rect 4920 15260 5296 15269
rect 4976 15258 5000 15260
rect 5056 15258 5080 15260
rect 5136 15258 5160 15260
rect 5216 15258 5240 15260
rect 4976 15206 4986 15258
rect 5230 15206 5240 15258
rect 4976 15204 5000 15206
rect 5056 15204 5080 15206
rect 5136 15204 5160 15206
rect 5216 15204 5240 15206
rect 4920 15195 5296 15204
rect 4920 14172 5296 14181
rect 4976 14170 5000 14172
rect 5056 14170 5080 14172
rect 5136 14170 5160 14172
rect 5216 14170 5240 14172
rect 4976 14118 4986 14170
rect 5230 14118 5240 14170
rect 4976 14116 5000 14118
rect 5056 14116 5080 14118
rect 5136 14116 5160 14118
rect 5216 14116 5240 14118
rect 4920 14107 5296 14116
rect 5460 13410 5488 16050
rect 5460 13382 5672 13410
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 4920 13084 5296 13093
rect 4976 13082 5000 13084
rect 5056 13082 5080 13084
rect 5136 13082 5160 13084
rect 5216 13082 5240 13084
rect 4976 13030 4986 13082
rect 5230 13030 5240 13082
rect 4976 13028 5000 13030
rect 5056 13028 5080 13030
rect 5136 13028 5160 13030
rect 5216 13028 5240 13030
rect 4920 13019 5296 13028
rect 5368 12850 5396 13126
rect 5552 12986 5580 13262
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 4528 12776 4580 12782
rect 4580 12724 4660 12730
rect 4528 12718 4660 12724
rect 4540 12702 4660 12718
rect 4180 12540 4556 12549
rect 4236 12538 4260 12540
rect 4316 12538 4340 12540
rect 4396 12538 4420 12540
rect 4476 12538 4500 12540
rect 4236 12486 4246 12538
rect 4490 12486 4500 12538
rect 4236 12484 4260 12486
rect 4316 12484 4340 12486
rect 4396 12484 4420 12486
rect 4476 12484 4500 12486
rect 4180 12475 4556 12484
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3804 10742 3832 11494
rect 4180 11452 4556 11461
rect 4236 11450 4260 11452
rect 4316 11450 4340 11452
rect 4396 11450 4420 11452
rect 4476 11450 4500 11452
rect 4236 11398 4246 11450
rect 4490 11398 4500 11450
rect 4236 11396 4260 11398
rect 4316 11396 4340 11398
rect 4396 11396 4420 11398
rect 4476 11396 4500 11398
rect 4180 11387 4556 11396
rect 4632 11354 4660 12702
rect 4724 12102 4752 12838
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5460 12442 5488 12854
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5552 12434 5580 12582
rect 5644 12434 5672 13382
rect 5552 12406 5672 12434
rect 5552 12322 5580 12406
rect 5368 12294 5580 12322
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4920 11996 5296 12005
rect 4976 11994 5000 11996
rect 5056 11994 5080 11996
rect 5136 11994 5160 11996
rect 5216 11994 5240 11996
rect 4976 11942 4986 11994
rect 5230 11942 5240 11994
rect 4976 11940 5000 11942
rect 5056 11940 5080 11942
rect 5136 11940 5160 11942
rect 5216 11940 5240 11942
rect 4920 11931 5296 11940
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 8906 2360 9318
rect 3344 8974 3372 10542
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3804 9382 3832 9522
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2792 8566 2820 8910
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 8090 2728 8434
rect 3804 8362 3832 9318
rect 3988 8430 4016 10610
rect 4080 10266 4108 10678
rect 4448 10470 4476 11290
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4540 10538 4568 11154
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4180 10364 4556 10373
rect 4236 10362 4260 10364
rect 4316 10362 4340 10364
rect 4396 10362 4420 10364
rect 4476 10362 4500 10364
rect 4236 10310 4246 10362
rect 4490 10310 4500 10362
rect 4236 10308 4260 10310
rect 4316 10308 4340 10310
rect 4396 10308 4420 10310
rect 4476 10308 4500 10310
rect 4180 10299 4556 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9450 4384 10066
rect 4632 10062 4660 11018
rect 4724 10810 4752 11086
rect 4816 10810 4844 11698
rect 4920 10908 5296 10917
rect 4976 10906 5000 10908
rect 5056 10906 5080 10908
rect 5136 10906 5160 10908
rect 5216 10906 5240 10908
rect 4976 10854 4986 10906
rect 5230 10854 5240 10906
rect 4976 10852 5000 10854
rect 5056 10852 5080 10854
rect 5136 10852 5160 10854
rect 5216 10852 5240 10854
rect 4920 10843 5296 10852
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4724 10062 4752 10746
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4816 10062 4844 10474
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10062 4936 10406
rect 5368 10062 5396 12294
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 10266 5488 12038
rect 5552 11898 5580 12106
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10810 5672 10950
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4180 9276 4556 9285
rect 4236 9274 4260 9276
rect 4316 9274 4340 9276
rect 4396 9274 4420 9276
rect 4476 9274 4500 9276
rect 4236 9222 4246 9274
rect 4490 9222 4500 9274
rect 4236 9220 4260 9222
rect 4316 9220 4340 9222
rect 4396 9220 4420 9222
rect 4476 9220 4500 9222
rect 4180 9211 4556 9220
rect 4724 9110 4752 9318
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4080 8634 4108 8774
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4632 8566 4660 8774
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4724 8498 4752 9046
rect 4816 8498 4844 9862
rect 4920 9820 5296 9829
rect 4976 9818 5000 9820
rect 5056 9818 5080 9820
rect 5136 9818 5160 9820
rect 5216 9818 5240 9820
rect 4976 9766 4986 9818
rect 5230 9766 5240 9818
rect 4976 9764 5000 9766
rect 5056 9764 5080 9766
rect 5136 9764 5160 9766
rect 5216 9764 5240 9766
rect 4920 9755 5296 9764
rect 4920 8732 5296 8741
rect 4976 8730 5000 8732
rect 5056 8730 5080 8732
rect 5136 8730 5160 8732
rect 5216 8730 5240 8732
rect 4976 8678 4986 8730
rect 5230 8678 5240 8730
rect 4976 8676 5000 8678
rect 5056 8676 5080 8678
rect 5136 8676 5160 8678
rect 5216 8676 5240 8678
rect 4920 8667 5296 8676
rect 5368 8498 5396 9998
rect 5736 9586 5764 20742
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5920 17610 5948 18022
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5816 15428 5868 15434
rect 5816 15370 5868 15376
rect 5828 15162 5856 15370
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 6012 12986 6040 13262
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6104 12434 6132 20402
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 20058 6408 20198
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6472 18630 6500 24670
rect 6564 18970 6592 27270
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 6644 25424 6696 25430
rect 6644 25366 6696 25372
rect 6656 24886 6684 25366
rect 7024 25242 7052 25638
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 6932 25214 7052 25242
rect 6644 24880 6696 24886
rect 6644 24822 6696 24828
rect 6840 23186 6868 25162
rect 6932 25158 6960 25214
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 7208 24750 7236 27406
rect 7392 25906 7420 28018
rect 7484 27606 7512 28562
rect 7656 28076 7708 28082
rect 7656 28018 7708 28024
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7392 25498 7420 25842
rect 7380 25492 7432 25498
rect 7380 25434 7432 25440
rect 7392 24886 7420 25434
rect 7484 25362 7512 27542
rect 7668 27470 7696 28018
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7760 27470 7788 27882
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7852 27538 7880 27814
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7656 27464 7708 27470
rect 7656 27406 7708 27412
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7380 24880 7432 24886
rect 7380 24822 7432 24828
rect 7668 24818 7696 27406
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7196 24744 7248 24750
rect 7196 24686 7248 24692
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6932 24410 6960 24550
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 6748 22778 6776 22918
rect 6736 22772 6788 22778
rect 6736 22714 6788 22720
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6656 21010 6684 21490
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6656 20602 6684 20946
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6840 20398 6868 23122
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20602 6960 20742
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 20058 6868 20334
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6564 18426 6592 18906
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6460 18148 6512 18154
rect 6460 18090 6512 18096
rect 6472 17134 6500 18090
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6564 17338 6592 17546
rect 6748 17338 6776 18362
rect 6840 18222 6868 18634
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6840 17218 6868 18158
rect 6748 17190 6868 17218
rect 7024 17218 7052 23258
rect 7208 22778 7236 24686
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7208 22094 7236 22714
rect 7668 22642 7696 24754
rect 7748 23044 7800 23050
rect 7748 22986 7800 22992
rect 7760 22778 7788 22986
rect 7748 22772 7800 22778
rect 7748 22714 7800 22720
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 22094 7696 22578
rect 7208 22066 7420 22094
rect 7392 22030 7420 22066
rect 7576 22066 7696 22094
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7392 21622 7420 21966
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7576 21554 7604 22066
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7116 20942 7144 21422
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7472 20868 7524 20874
rect 7472 20810 7524 20816
rect 7484 20602 7512 20810
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7576 19514 7604 21490
rect 7668 20466 7696 21830
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 8036 18290 8064 30194
rect 8484 29640 8536 29646
rect 8484 29582 8536 29588
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 8312 29306 8340 29446
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8496 28762 8524 29582
rect 8484 28756 8536 28762
rect 8484 28698 8536 28704
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8312 28218 8340 28358
rect 8404 28218 8432 28562
rect 8484 28484 8536 28490
rect 8484 28426 8536 28432
rect 8300 28212 8352 28218
rect 8300 28154 8352 28160
rect 8392 28212 8444 28218
rect 8392 28154 8444 28160
rect 8116 25900 8168 25906
rect 8116 25842 8168 25848
rect 8128 25498 8156 25842
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 8128 23730 8156 24822
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 23866 8432 24006
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8128 23118 8156 23666
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8128 21010 8156 22034
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21690 8248 21830
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8312 19854 8340 21286
rect 8404 21146 8432 21286
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8496 20890 8524 28426
rect 8588 28082 8616 30534
rect 8956 30394 8984 30534
rect 8944 30388 8996 30394
rect 8944 30330 8996 30336
rect 9140 28966 9168 30534
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9404 29504 9456 29510
rect 9404 29446 9456 29452
rect 9324 29306 9352 29446
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9416 28558 9444 29446
rect 9692 29102 9720 30738
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 10060 29646 10088 30670
rect 10428 30190 10456 30806
rect 10980 30734 11008 31078
rect 12912 30938 12940 31214
rect 14556 31204 14608 31210
rect 14556 31146 14608 31152
rect 16948 31204 17000 31210
rect 16948 31146 17000 31152
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 11888 30660 11940 30666
rect 11888 30602 11940 30608
rect 12808 30660 12860 30666
rect 12808 30602 12860 30608
rect 10920 30492 11296 30501
rect 10976 30490 11000 30492
rect 11056 30490 11080 30492
rect 11136 30490 11160 30492
rect 11216 30490 11240 30492
rect 10976 30438 10986 30490
rect 11230 30438 11240 30490
rect 10976 30436 11000 30438
rect 11056 30436 11080 30438
rect 11136 30436 11160 30438
rect 11216 30436 11240 30438
rect 10920 30427 11296 30436
rect 11900 30326 11928 30602
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12084 30410 12112 30534
rect 12084 30394 12296 30410
rect 12084 30388 12308 30394
rect 12084 30382 12256 30388
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 10416 30184 10468 30190
rect 10416 30126 10468 30132
rect 10784 30184 10836 30190
rect 10784 30126 10836 30132
rect 10180 29948 10556 29957
rect 10236 29946 10260 29948
rect 10316 29946 10340 29948
rect 10396 29946 10420 29948
rect 10476 29946 10500 29948
rect 10236 29894 10246 29946
rect 10490 29894 10500 29946
rect 10236 29892 10260 29894
rect 10316 29892 10340 29894
rect 10396 29892 10420 29894
rect 10476 29892 10500 29894
rect 10180 29883 10556 29892
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 8772 27674 8800 28018
rect 9140 27674 9168 28018
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 9588 26376 9640 26382
rect 9692 26364 9720 29038
rect 10180 28860 10556 28869
rect 10236 28858 10260 28860
rect 10316 28858 10340 28860
rect 10396 28858 10420 28860
rect 10476 28858 10500 28860
rect 10236 28806 10246 28858
rect 10490 28806 10500 28858
rect 10236 28804 10260 28806
rect 10316 28804 10340 28806
rect 10396 28804 10420 28806
rect 10476 28804 10500 28806
rect 10180 28795 10556 28804
rect 10612 28762 10640 29106
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 9956 28620 10008 28626
rect 9956 28562 10008 28568
rect 9640 26336 9720 26364
rect 9588 26318 9640 26324
rect 8588 26042 8616 26318
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23866 8616 24142
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8864 22094 8892 25638
rect 9324 25498 9352 25638
rect 9600 25498 9628 26318
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9324 24954 9352 25230
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9692 24886 9720 25842
rect 9968 25838 9996 28562
rect 10704 27946 10732 29446
rect 10692 27940 10744 27946
rect 10692 27882 10744 27888
rect 10180 27772 10556 27781
rect 10236 27770 10260 27772
rect 10316 27770 10340 27772
rect 10396 27770 10420 27772
rect 10476 27770 10500 27772
rect 10236 27718 10246 27770
rect 10490 27718 10500 27770
rect 10236 27716 10260 27718
rect 10316 27716 10340 27718
rect 10396 27716 10420 27718
rect 10476 27716 10500 27718
rect 10180 27707 10556 27716
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 10692 26784 10744 26790
rect 10692 26726 10744 26732
rect 10060 26042 10088 26726
rect 10180 26684 10556 26693
rect 10236 26682 10260 26684
rect 10316 26682 10340 26684
rect 10396 26682 10420 26684
rect 10476 26682 10500 26684
rect 10236 26630 10246 26682
rect 10490 26630 10500 26682
rect 10236 26628 10260 26630
rect 10316 26628 10340 26630
rect 10396 26628 10420 26630
rect 10476 26628 10500 26630
rect 10180 26619 10556 26628
rect 10704 26518 10732 26726
rect 10692 26512 10744 26518
rect 10692 26454 10744 26460
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10428 26042 10456 26182
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 9956 25832 10008 25838
rect 9876 25792 9956 25820
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9692 24750 9720 24822
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 9692 23866 9720 24006
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9876 23662 9904 25792
rect 9956 25774 10008 25780
rect 10520 25770 10548 26318
rect 10600 25832 10652 25838
rect 10796 25820 10824 30126
rect 11532 30122 11560 30194
rect 11520 30116 11572 30122
rect 11520 30058 11572 30064
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 10920 29404 11296 29413
rect 10976 29402 11000 29404
rect 11056 29402 11080 29404
rect 11136 29402 11160 29404
rect 11216 29402 11240 29404
rect 10976 29350 10986 29402
rect 11230 29350 11240 29402
rect 10976 29348 11000 29350
rect 11056 29348 11080 29350
rect 11136 29348 11160 29350
rect 11216 29348 11240 29350
rect 10920 29339 11296 29348
rect 11348 28694 11376 29582
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11716 29306 11744 29446
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11992 29102 12020 29786
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11336 28688 11388 28694
rect 11336 28630 11388 28636
rect 10920 28316 11296 28325
rect 10976 28314 11000 28316
rect 11056 28314 11080 28316
rect 11136 28314 11160 28316
rect 11216 28314 11240 28316
rect 10976 28262 10986 28314
rect 11230 28262 11240 28314
rect 10976 28260 11000 28262
rect 11056 28260 11080 28262
rect 11136 28260 11160 28262
rect 11216 28260 11240 28262
rect 10920 28251 11296 28260
rect 11152 27872 11204 27878
rect 11152 27814 11204 27820
rect 11164 27418 11192 27814
rect 11348 27554 11376 28630
rect 11532 28558 11560 28902
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 11624 27878 11652 28902
rect 11992 28490 12020 29038
rect 12084 28558 12112 30382
rect 12256 30330 12308 30336
rect 12360 30258 12388 30534
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 12820 30054 12848 30602
rect 12808 30048 12860 30054
rect 12808 29990 12860 29996
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12256 29572 12308 29578
rect 12256 29514 12308 29520
rect 12164 29096 12216 29102
rect 12164 29038 12216 29044
rect 12176 28626 12204 29038
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 12164 28484 12216 28490
rect 12268 28472 12296 29514
rect 12360 29102 12388 29582
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12544 29306 12572 29446
rect 12532 29300 12584 29306
rect 12532 29242 12584 29248
rect 12912 29170 12940 30874
rect 14004 30728 14056 30734
rect 14004 30670 14056 30676
rect 14016 30394 14044 30670
rect 14004 30388 14056 30394
rect 14004 30330 14056 30336
rect 14568 30190 14596 31146
rect 16180 31036 16556 31045
rect 16236 31034 16260 31036
rect 16316 31034 16340 31036
rect 16396 31034 16420 31036
rect 16476 31034 16500 31036
rect 16236 30982 16246 31034
rect 16490 30982 16500 31034
rect 16236 30980 16260 30982
rect 16316 30980 16340 30982
rect 16396 30980 16420 30982
rect 16476 30980 16500 30982
rect 16180 30971 16556 30980
rect 16960 30938 16988 31146
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17604 30938 17632 31078
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14660 29646 14688 30670
rect 15016 30592 15068 30598
rect 15016 30534 15068 30540
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14660 29306 14688 29582
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 14936 29306 14964 29514
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14924 29300 14976 29306
rect 14924 29242 14976 29248
rect 12900 29164 12952 29170
rect 12900 29106 12952 29112
rect 13176 29164 13228 29170
rect 13176 29106 13228 29112
rect 12348 29096 12400 29102
rect 12348 29038 12400 29044
rect 12360 28558 12388 29038
rect 13084 28960 13136 28966
rect 13084 28902 13136 28908
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12216 28444 12296 28472
rect 12164 28426 12216 28432
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11348 27526 11468 27554
rect 11164 27390 11376 27418
rect 10920 27228 11296 27237
rect 10976 27226 11000 27228
rect 11056 27226 11080 27228
rect 11136 27226 11160 27228
rect 11216 27226 11240 27228
rect 10976 27174 10986 27226
rect 11230 27174 11240 27226
rect 10976 27172 11000 27174
rect 11056 27172 11080 27174
rect 11136 27172 11160 27174
rect 11216 27172 11240 27174
rect 10920 27163 11296 27172
rect 10920 26140 11296 26149
rect 10976 26138 11000 26140
rect 11056 26138 11080 26140
rect 11136 26138 11160 26140
rect 11216 26138 11240 26140
rect 10976 26086 10986 26138
rect 11230 26086 11240 26138
rect 10976 26084 11000 26086
rect 11056 26084 11080 26086
rect 11136 26084 11160 26086
rect 11216 26084 11240 26086
rect 10920 26075 11296 26084
rect 10652 25792 10824 25820
rect 10600 25774 10652 25780
rect 10508 25764 10560 25770
rect 10508 25706 10560 25712
rect 10180 25596 10556 25605
rect 10236 25594 10260 25596
rect 10316 25594 10340 25596
rect 10396 25594 10420 25596
rect 10476 25594 10500 25596
rect 10236 25542 10246 25594
rect 10490 25542 10500 25594
rect 10236 25540 10260 25542
rect 10316 25540 10340 25542
rect 10396 25540 10420 25542
rect 10476 25540 10500 25542
rect 10180 25531 10556 25540
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9968 24954 9996 25094
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 10140 24744 10192 24750
rect 10060 24692 10140 24698
rect 10060 24686 10192 24692
rect 10060 24670 10180 24686
rect 9956 23724 10008 23730
rect 9956 23666 10008 23672
rect 9864 23656 9916 23662
rect 9692 23604 9864 23610
rect 9692 23598 9916 23604
rect 9692 23582 9904 23598
rect 9220 23520 9272 23526
rect 9220 23462 9272 23468
rect 9232 23186 9260 23462
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8956 22778 8984 22918
rect 8944 22772 8996 22778
rect 8944 22714 8996 22720
rect 8864 22066 8984 22094
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8404 20862 8524 20890
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8404 18358 8432 20862
rect 8772 20806 8800 21422
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8496 20466 8524 20742
rect 8772 20466 8800 20742
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7024 17190 7144 17218
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15706 6408 15846
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6656 15162 6684 16186
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6748 14890 6776 17190
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16726 6868 17070
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6840 16046 6868 16662
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6736 14884 6788 14890
rect 6736 14826 6788 14832
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 5920 12406 6132 12434
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8634 5672 8774
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 3896 7886 3924 8230
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 4080 6186 4108 8366
rect 4180 8188 4556 8197
rect 4236 8186 4260 8188
rect 4316 8186 4340 8188
rect 4396 8186 4420 8188
rect 4476 8186 4500 8188
rect 4236 8134 4246 8186
rect 4490 8134 4500 8186
rect 4236 8132 4260 8134
rect 4316 8132 4340 8134
rect 4396 8132 4420 8134
rect 4476 8132 4500 8134
rect 4180 8123 4556 8132
rect 4920 7644 5296 7653
rect 4976 7642 5000 7644
rect 5056 7642 5080 7644
rect 5136 7642 5160 7644
rect 5216 7642 5240 7644
rect 4976 7590 4986 7642
rect 5230 7590 5240 7642
rect 4976 7588 5000 7590
rect 5056 7588 5080 7590
rect 5136 7588 5160 7590
rect 5216 7588 5240 7590
rect 4920 7579 5296 7588
rect 4180 7100 4556 7109
rect 4236 7098 4260 7100
rect 4316 7098 4340 7100
rect 4396 7098 4420 7100
rect 4476 7098 4500 7100
rect 4236 7046 4246 7098
rect 4490 7046 4500 7098
rect 4236 7044 4260 7046
rect 4316 7044 4340 7046
rect 4396 7044 4420 7046
rect 4476 7044 4500 7046
rect 4180 7035 4556 7044
rect 5920 6798 5948 12406
rect 6196 12374 6224 13194
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6472 12714 6500 13126
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9586 6408 9862
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6012 9042 6040 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6012 8634 6040 8978
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 4920 6556 5296 6565
rect 4976 6554 5000 6556
rect 5056 6554 5080 6556
rect 5136 6554 5160 6556
rect 5216 6554 5240 6556
rect 4976 6502 4986 6554
rect 5230 6502 5240 6554
rect 4976 6500 5000 6502
rect 5056 6500 5080 6502
rect 5136 6500 5160 6502
rect 5216 6500 5240 6502
rect 4920 6491 5296 6500
rect 5920 6458 5948 6734
rect 6012 6458 6040 8570
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 4080 5574 4108 6122
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 4180 6012 4556 6021
rect 4236 6010 4260 6012
rect 4316 6010 4340 6012
rect 4396 6010 4420 6012
rect 4476 6010 4500 6012
rect 4236 5958 4246 6010
rect 4490 5958 4500 6010
rect 4236 5956 4260 5958
rect 4316 5956 4340 5958
rect 4396 5956 4420 5958
rect 4476 5956 4500 5958
rect 4180 5947 4556 5956
rect 5368 5914 5396 6054
rect 6012 5914 6040 6394
rect 6196 6254 6224 9114
rect 6564 8974 6592 9318
rect 6656 9178 6684 12718
rect 6748 12434 6776 14826
rect 6840 12782 6868 15982
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6748 12406 6868 12434
rect 6840 12306 6868 12406
rect 7024 12306 7052 12854
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6840 9518 6868 12242
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6840 6866 6868 9454
rect 6932 7886 6960 10542
rect 7116 9654 7144 17190
rect 8036 17105 8064 18226
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17542 8156 18158
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 17270 8156 17478
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8220 17202 8248 17750
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8312 17338 8340 17478
rect 8404 17338 8432 18294
rect 8772 18222 8800 20402
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8022 17096 8078 17105
rect 8022 17031 8078 17040
rect 8036 16794 8064 17031
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7300 15026 7328 15914
rect 7852 15706 7880 15982
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7760 15026 7788 15302
rect 7852 15162 7880 15642
rect 7944 15570 7972 15982
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 8220 15094 8248 17138
rect 8404 16250 8432 17274
rect 8772 17202 8800 18158
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 8220 14890 8248 15030
rect 8496 15026 8524 17138
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 8208 14884 8260 14890
rect 8208 14826 8260 14832
rect 7300 13326 7328 14826
rect 8496 13802 8524 14962
rect 8956 14074 8984 22066
rect 9312 22024 9364 22030
rect 9692 21978 9720 23582
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9784 23186 9812 23462
rect 9968 23322 9996 23666
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9784 22234 9812 23122
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9312 21966 9364 21972
rect 9324 21146 9352 21966
rect 9600 21950 9720 21978
rect 9600 21434 9628 21950
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9692 21554 9720 21830
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9600 21406 9720 21434
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9692 21049 9720 21406
rect 9678 21040 9734 21049
rect 9678 20975 9734 20984
rect 9784 20942 9812 21830
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9692 20602 9720 20878
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9140 18426 9168 18566
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9324 17882 9352 18702
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 17649 9628 17682
rect 9586 17640 9642 17649
rect 9586 17575 9642 17584
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9140 16794 9168 17206
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9600 16658 9628 17206
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9600 15162 9628 15370
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 8944 14068 8996 14074
rect 8996 14028 9076 14056
rect 8944 14010 8996 14016
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 7748 13524 7800 13530
rect 7852 13512 7880 13738
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 7800 13484 7880 13512
rect 7748 13466 7800 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7208 12986 7236 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7208 9722 7236 9862
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7300 9654 7328 13262
rect 7392 12918 7420 13262
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7116 8974 7144 9590
rect 7760 9586 7788 9998
rect 7852 9586 7880 13484
rect 8680 13394 8708 13670
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 7944 12442 7972 12854
rect 8220 12442 8248 13194
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7944 11218 7972 12378
rect 8864 12238 8892 12582
rect 8956 12374 8984 13126
rect 9048 12986 9076 14028
rect 9692 13954 9720 17750
rect 9784 17746 9812 18702
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9600 13926 9720 13954
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13326 9168 13670
rect 9600 13462 9628 13926
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9692 13530 9720 13806
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 12434 9444 12922
rect 9416 12406 9628 12434
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 9600 11762 9628 12406
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11762 9720 12038
rect 9784 11762 9812 15982
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8772 11150 8800 11494
rect 9600 11150 9628 11698
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9692 10810 9720 11562
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9876 10010 9904 23054
rect 10060 21690 10088 24670
rect 10180 24508 10556 24517
rect 10236 24506 10260 24508
rect 10316 24506 10340 24508
rect 10396 24506 10420 24508
rect 10476 24506 10500 24508
rect 10236 24454 10246 24506
rect 10490 24454 10500 24506
rect 10236 24452 10260 24454
rect 10316 24452 10340 24454
rect 10396 24452 10420 24454
rect 10476 24452 10500 24454
rect 10180 24443 10556 24452
rect 10612 23526 10640 25774
rect 10920 25052 11296 25061
rect 10976 25050 11000 25052
rect 11056 25050 11080 25052
rect 11136 25050 11160 25052
rect 11216 25050 11240 25052
rect 10976 24998 10986 25050
rect 11230 24998 11240 25050
rect 10976 24996 11000 24998
rect 11056 24996 11080 24998
rect 11136 24996 11160 24998
rect 11216 24996 11240 24998
rect 10920 24987 11296 24996
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10704 23633 10732 24754
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10690 23624 10746 23633
rect 10796 23594 10824 24142
rect 10920 23964 11296 23973
rect 10976 23962 11000 23964
rect 11056 23962 11080 23964
rect 11136 23962 11160 23964
rect 11216 23962 11240 23964
rect 10976 23910 10986 23962
rect 11230 23910 11240 23962
rect 10976 23908 11000 23910
rect 11056 23908 11080 23910
rect 11136 23908 11160 23910
rect 11216 23908 11240 23910
rect 10920 23899 11296 23908
rect 10690 23559 10746 23568
rect 10784 23588 10836 23594
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10180 23420 10556 23429
rect 10236 23418 10260 23420
rect 10316 23418 10340 23420
rect 10396 23418 10420 23420
rect 10476 23418 10500 23420
rect 10236 23366 10246 23418
rect 10490 23366 10500 23418
rect 10236 23364 10260 23366
rect 10316 23364 10340 23366
rect 10396 23364 10420 23366
rect 10476 23364 10500 23366
rect 10180 23355 10556 23364
rect 10232 23112 10284 23118
rect 10230 23080 10232 23089
rect 10600 23112 10652 23118
rect 10284 23080 10286 23089
rect 10600 23054 10652 23060
rect 10230 23015 10286 23024
rect 10180 22332 10556 22341
rect 10236 22330 10260 22332
rect 10316 22330 10340 22332
rect 10396 22330 10420 22332
rect 10476 22330 10500 22332
rect 10236 22278 10246 22330
rect 10490 22278 10500 22330
rect 10236 22276 10260 22278
rect 10316 22276 10340 22278
rect 10396 22276 10420 22278
rect 10476 22276 10500 22278
rect 10180 22267 10556 22276
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 19854 9996 21286
rect 10060 21010 10088 21626
rect 10180 21244 10556 21253
rect 10236 21242 10260 21244
rect 10316 21242 10340 21244
rect 10396 21242 10420 21244
rect 10476 21242 10500 21244
rect 10236 21190 10246 21242
rect 10490 21190 10500 21242
rect 10236 21188 10260 21190
rect 10316 21188 10340 21190
rect 10396 21188 10420 21190
rect 10476 21188 10500 21190
rect 10180 21179 10556 21188
rect 10322 21040 10378 21049
rect 10048 21004 10100 21010
rect 10322 20975 10378 20984
rect 10048 20946 10100 20952
rect 10336 20398 10364 20975
rect 10612 20913 10640 23054
rect 10704 21554 10732 23559
rect 10784 23530 10836 23536
rect 10796 23118 10824 23530
rect 10876 23316 10928 23322
rect 10876 23258 10928 23264
rect 10888 23118 10916 23258
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10920 22876 11296 22885
rect 10976 22874 11000 22876
rect 11056 22874 11080 22876
rect 11136 22874 11160 22876
rect 11216 22874 11240 22876
rect 10976 22822 10986 22874
rect 11230 22822 11240 22874
rect 10976 22820 11000 22822
rect 11056 22820 11080 22822
rect 11136 22820 11160 22822
rect 11216 22820 11240 22822
rect 10920 22811 11296 22820
rect 10784 22160 10836 22166
rect 10784 22102 10836 22108
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10704 20942 10732 21490
rect 10692 20936 10744 20942
rect 10598 20904 10654 20913
rect 10692 20878 10744 20884
rect 10598 20839 10654 20848
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10180 20156 10556 20165
rect 10236 20154 10260 20156
rect 10316 20154 10340 20156
rect 10396 20154 10420 20156
rect 10476 20154 10500 20156
rect 10236 20102 10246 20154
rect 10490 20102 10500 20154
rect 10236 20100 10260 20102
rect 10316 20100 10340 20102
rect 10396 20100 10420 20102
rect 10476 20100 10500 20102
rect 10180 20091 10556 20100
rect 10612 19854 10640 20839
rect 10796 20584 10824 22102
rect 10920 21788 11296 21797
rect 10976 21786 11000 21788
rect 11056 21786 11080 21788
rect 11136 21786 11160 21788
rect 11216 21786 11240 21788
rect 10976 21734 10986 21786
rect 11230 21734 11240 21786
rect 10976 21732 11000 21734
rect 11056 21732 11080 21734
rect 11136 21732 11160 21734
rect 11216 21732 11240 21734
rect 10920 21723 11296 21732
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11072 20874 11100 21422
rect 11060 20868 11112 20874
rect 11060 20810 11112 20816
rect 10920 20700 11296 20709
rect 10976 20698 11000 20700
rect 11056 20698 11080 20700
rect 11136 20698 11160 20700
rect 11216 20698 11240 20700
rect 10976 20646 10986 20698
rect 11230 20646 11240 20698
rect 10976 20644 11000 20646
rect 11056 20644 11080 20646
rect 11136 20644 11160 20646
rect 11216 20644 11240 20646
rect 10920 20635 11296 20644
rect 10796 20556 10916 20584
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10796 19990 10824 20402
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10888 19854 10916 20556
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 11348 19666 11376 27390
rect 11440 26586 11468 27526
rect 11980 27464 12032 27470
rect 11980 27406 12032 27412
rect 11992 27130 12020 27406
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 20942 11468 24550
rect 11532 23322 11560 26318
rect 12176 26314 12204 28426
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 11704 26240 11756 26246
rect 11704 26182 11756 26188
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11624 24818 11652 25298
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11716 24206 11744 26182
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11532 22166 11560 23258
rect 11704 23180 11756 23186
rect 11808 23168 11836 26250
rect 12360 25838 12388 27406
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12452 25906 12480 26318
rect 12900 26240 12952 26246
rect 12900 26182 12952 26188
rect 12912 25974 12940 26182
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11992 24614 12020 25638
rect 12360 25498 12388 25774
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24954 12388 25162
rect 12452 24954 12480 25842
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12544 25158 12572 25774
rect 13096 25702 13124 28902
rect 13188 28762 13216 29106
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 14476 28626 14504 29242
rect 13176 28620 13228 28626
rect 13176 28562 13228 28568
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 13188 27062 13216 28562
rect 15028 28558 15056 30534
rect 15580 30394 15608 30534
rect 16920 30492 17296 30501
rect 16976 30490 17000 30492
rect 17056 30490 17080 30492
rect 17136 30490 17160 30492
rect 17216 30490 17240 30492
rect 16976 30438 16986 30490
rect 17230 30438 17240 30490
rect 16976 30436 17000 30438
rect 17056 30436 17080 30438
rect 17136 30436 17160 30438
rect 17216 30436 17240 30438
rect 16920 30427 17296 30436
rect 15568 30388 15620 30394
rect 15568 30330 15620 30336
rect 17328 30258 17356 30670
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17420 30394 17448 30534
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 16180 29948 16556 29957
rect 16236 29946 16260 29948
rect 16316 29946 16340 29948
rect 16396 29946 16420 29948
rect 16476 29946 16500 29948
rect 16236 29894 16246 29946
rect 16490 29894 16500 29946
rect 16236 29892 16260 29894
rect 16316 29892 16340 29894
rect 16396 29892 16420 29894
rect 16476 29892 16500 29894
rect 16180 29883 16556 29892
rect 15292 29844 15344 29850
rect 15292 29786 15344 29792
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15108 28960 15160 28966
rect 15108 28902 15160 28908
rect 15120 28558 15148 28902
rect 15212 28558 15240 29446
rect 15304 29306 15332 29786
rect 17328 29646 17356 30194
rect 17972 30054 18000 31214
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 17316 29640 17368 29646
rect 17316 29582 17368 29588
rect 15384 29572 15436 29578
rect 15384 29514 15436 29520
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 14556 28416 14608 28422
rect 14556 28358 14608 28364
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13176 27056 13228 27062
rect 13176 26998 13228 27004
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12544 24886 12572 25094
rect 12532 24880 12584 24886
rect 12532 24822 12584 24828
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 12084 24410 12112 24550
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 11756 23140 11836 23168
rect 11704 23122 11756 23128
rect 11612 23044 11664 23050
rect 11612 22986 11664 22992
rect 11624 22778 11652 22986
rect 11612 22772 11664 22778
rect 11612 22714 11664 22720
rect 11900 22710 11928 23190
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 12084 22522 12112 22918
rect 11900 22494 12112 22522
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11532 21978 11560 22102
rect 11532 21950 11836 21978
rect 11808 21894 11836 21950
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11624 21350 11652 21830
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11624 20942 11652 21286
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11440 20058 11468 20742
rect 11716 20466 11744 21422
rect 11900 21298 11928 22494
rect 12176 22386 12204 24754
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23202 12296 24006
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12268 23174 12388 23202
rect 12452 23186 12480 23462
rect 12544 23186 12572 24822
rect 13464 24682 13492 25094
rect 13556 24818 13584 27950
rect 13648 27674 13676 28086
rect 13728 28076 13780 28082
rect 13728 28018 13780 28024
rect 13636 27668 13688 27674
rect 13636 27610 13688 27616
rect 13740 27606 13768 28018
rect 13728 27600 13780 27606
rect 13728 27542 13780 27548
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13648 26518 13676 26726
rect 13636 26512 13688 26518
rect 13636 26454 13688 26460
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13372 24410 13400 24550
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13464 23730 13492 23802
rect 13556 23730 13584 24754
rect 13740 24682 13768 27542
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 27130 14136 27270
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24954 14136 25094
rect 14096 24948 14148 24954
rect 14096 24890 14148 24896
rect 14568 24750 14596 28358
rect 15200 26512 15252 26518
rect 15200 26454 15252 26460
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14660 26042 14688 26318
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14660 24954 14688 25978
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14648 24948 14700 24954
rect 14648 24890 14700 24896
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 13728 24676 13780 24682
rect 13728 24618 13780 24624
rect 13740 24070 13768 24618
rect 14372 24608 14424 24614
rect 14372 24550 14424 24556
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13740 23866 13768 24006
rect 13832 23866 13860 24074
rect 14384 23866 14412 24550
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12268 22778 12296 23054
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 11992 22358 12204 22386
rect 11992 21962 12020 22358
rect 12360 22094 12388 23174
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12624 23112 12676 23118
rect 12622 23080 12624 23089
rect 12676 23080 12678 23089
rect 12622 23015 12678 23024
rect 12820 22094 12848 23666
rect 14568 23662 14596 24686
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13464 22642 13492 23530
rect 13924 23322 13952 23598
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14108 22778 14136 22918
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12912 22166 12940 22442
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12084 22066 12388 22094
rect 12728 22066 12848 22094
rect 13268 22092 13320 22098
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11808 21270 11928 21298
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11348 19638 11560 19666
rect 10920 19612 11296 19621
rect 10976 19610 11000 19612
rect 11056 19610 11080 19612
rect 11136 19610 11160 19612
rect 11216 19610 11240 19612
rect 10976 19558 10986 19610
rect 11230 19558 11240 19610
rect 10976 19556 11000 19558
rect 11056 19556 11080 19558
rect 11136 19556 11160 19558
rect 11216 19556 11240 19558
rect 10920 19547 11296 19556
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9968 17678 9996 18090
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10060 17134 10088 19110
rect 10180 19068 10556 19077
rect 10236 19066 10260 19068
rect 10316 19066 10340 19068
rect 10396 19066 10420 19068
rect 10476 19066 10500 19068
rect 10236 19014 10246 19066
rect 10490 19014 10500 19066
rect 10236 19012 10260 19014
rect 10316 19012 10340 19014
rect 10396 19012 10420 19014
rect 10476 19012 10500 19014
rect 10180 19003 10556 19012
rect 10920 18524 11296 18533
rect 10976 18522 11000 18524
rect 11056 18522 11080 18524
rect 11136 18522 11160 18524
rect 11216 18522 11240 18524
rect 10976 18470 10986 18522
rect 11230 18470 11240 18522
rect 10976 18468 11000 18470
rect 11056 18468 11080 18470
rect 11136 18468 11160 18470
rect 11216 18468 11240 18470
rect 10920 18459 11296 18468
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10180 17980 10556 17989
rect 10236 17978 10260 17980
rect 10316 17978 10340 17980
rect 10396 17978 10420 17980
rect 10476 17978 10500 17980
rect 10236 17926 10246 17978
rect 10490 17926 10500 17978
rect 10236 17924 10260 17926
rect 10316 17924 10340 17926
rect 10396 17924 10420 17926
rect 10476 17924 10500 17926
rect 10180 17915 10556 17924
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 10152 17338 10180 17478
rect 10428 17338 10456 17478
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10612 17270 10640 18158
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 10920 17436 11296 17445
rect 10976 17434 11000 17436
rect 11056 17434 11080 17436
rect 11136 17434 11160 17436
rect 11216 17434 11240 17436
rect 10976 17382 10986 17434
rect 11230 17382 11240 17434
rect 10976 17380 11000 17382
rect 11056 17380 11080 17382
rect 11136 17380 11160 17382
rect 11216 17380 11240 17382
rect 10920 17371 11296 17380
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10874 17232 10930 17241
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10180 16892 10556 16901
rect 10236 16890 10260 16892
rect 10316 16890 10340 16892
rect 10396 16890 10420 16892
rect 10476 16890 10500 16892
rect 10236 16838 10246 16890
rect 10490 16838 10500 16890
rect 10236 16836 10260 16838
rect 10316 16836 10340 16838
rect 10396 16836 10420 16838
rect 10476 16836 10500 16838
rect 10180 16827 10556 16836
rect 10612 16674 10640 17206
rect 10874 17167 10930 17176
rect 10888 17134 10916 17167
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 10888 16810 10916 17070
rect 10336 16646 10640 16674
rect 10704 16782 10916 16810
rect 11164 16794 11192 17070
rect 11152 16788 11204 16794
rect 10336 16250 10364 16646
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10180 15804 10556 15813
rect 10236 15802 10260 15804
rect 10316 15802 10340 15804
rect 10396 15802 10420 15804
rect 10476 15802 10500 15804
rect 10236 15750 10246 15802
rect 10490 15750 10500 15802
rect 10236 15748 10260 15750
rect 10316 15748 10340 15750
rect 10396 15748 10420 15750
rect 10476 15748 10500 15750
rect 10180 15739 10556 15748
rect 10704 15586 10732 16782
rect 11152 16730 11204 16736
rect 11348 16538 11376 17478
rect 11426 17368 11482 17377
rect 11426 17303 11482 17312
rect 11440 17202 11468 17303
rect 11532 17202 11560 19638
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11624 17678 11652 18226
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17338 11652 17478
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 11256 16510 11376 16538
rect 10520 15558 10732 15586
rect 10796 15570 10824 16458
rect 11152 16448 11204 16454
rect 11256 16436 11284 16510
rect 11204 16408 11284 16436
rect 11336 16448 11388 16454
rect 11152 16390 11204 16396
rect 11336 16390 11388 16396
rect 10920 16348 11296 16357
rect 10976 16346 11000 16348
rect 11056 16346 11080 16348
rect 11136 16346 11160 16348
rect 11216 16346 11240 16348
rect 10976 16294 10986 16346
rect 11230 16294 11240 16346
rect 10976 16292 11000 16294
rect 11056 16292 11080 16294
rect 11136 16292 11160 16294
rect 11216 16292 11240 16294
rect 10920 16283 11296 16292
rect 11348 16250 11376 16390
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10980 15706 11008 16118
rect 11440 16046 11468 16594
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11532 15892 11560 16662
rect 11348 15864 11560 15892
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10784 15564 10836 15570
rect 10520 14906 10548 15558
rect 10784 15506 10836 15512
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 15450 10916 15506
rect 10796 15422 10916 15450
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15162 10732 15302
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10520 14878 10732 14906
rect 10180 14716 10556 14725
rect 10236 14714 10260 14716
rect 10316 14714 10340 14716
rect 10396 14714 10420 14716
rect 10476 14714 10500 14716
rect 10236 14662 10246 14714
rect 10490 14662 10500 14714
rect 10236 14660 10260 14662
rect 10316 14660 10340 14662
rect 10396 14660 10420 14662
rect 10476 14660 10500 14662
rect 10180 14651 10556 14660
rect 10180 13628 10556 13637
rect 10236 13626 10260 13628
rect 10316 13626 10340 13628
rect 10396 13626 10420 13628
rect 10476 13626 10500 13628
rect 10236 13574 10246 13626
rect 10490 13574 10500 13626
rect 10236 13572 10260 13574
rect 10316 13572 10340 13574
rect 10396 13572 10420 13574
rect 10476 13572 10500 13574
rect 10180 13563 10556 13572
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 13274 9996 13330
rect 10600 13320 10652 13326
rect 9968 13246 10088 13274
rect 10600 13262 10652 13268
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9968 12986 9996 13126
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11286 9996 11494
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9784 9982 9904 10010
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 9784 9602 9812 9982
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9722 9904 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7024 6798 7052 8230
rect 7116 8090 7144 8910
rect 7576 8634 7604 9522
rect 7760 9178 7788 9522
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8634 7880 8774
rect 7944 8634 7972 8910
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6254 6316 6598
rect 7944 6458 7972 6802
rect 8312 6798 8340 9590
rect 8484 9580 8536 9586
rect 9784 9574 9904 9602
rect 8484 9522 8536 9528
rect 8496 6798 8524 9522
rect 9876 9518 9904 9574
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9324 9178 9352 9318
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8498 8708 8842
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8498 8892 8774
rect 9232 8634 9260 8910
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 8668 8492 8720 8498
rect 8852 8492 8904 8498
rect 8720 8452 8800 8480
rect 8668 8434 8720 8440
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6458 8064 6598
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6380 5914 6408 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 8036 5710 8064 6394
rect 8128 5914 8156 6734
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 6458 8708 6598
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 4068 5568 4120 5574
rect 1398 5536 1454 5545
rect 4068 5510 4120 5516
rect 1398 5471 1454 5480
rect 4920 5468 5296 5477
rect 4976 5466 5000 5468
rect 5056 5466 5080 5468
rect 5136 5466 5160 5468
rect 5216 5466 5240 5468
rect 4976 5414 4986 5466
rect 5230 5414 5240 5466
rect 4976 5412 5000 5414
rect 5056 5412 5080 5414
rect 5136 5412 5160 5414
rect 5216 5412 5240 5414
rect 4920 5403 5296 5412
rect 8772 5234 8800 8452
rect 8852 8434 8904 8440
rect 9876 7886 9904 9454
rect 9968 8906 9996 9998
rect 10060 9518 10088 13246
rect 10506 12880 10562 12889
rect 10506 12815 10508 12824
rect 10560 12815 10562 12824
rect 10508 12786 10560 12792
rect 10180 12540 10556 12549
rect 10236 12538 10260 12540
rect 10316 12538 10340 12540
rect 10396 12538 10420 12540
rect 10476 12538 10500 12540
rect 10236 12486 10246 12538
rect 10490 12486 10500 12538
rect 10236 12484 10260 12486
rect 10316 12484 10340 12486
rect 10396 12484 10420 12486
rect 10476 12484 10500 12486
rect 10180 12475 10556 12484
rect 10612 12442 10640 13262
rect 10704 12986 10732 14878
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10796 12866 10824 15422
rect 10980 15366 11008 15642
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10920 15260 11296 15269
rect 10976 15258 11000 15260
rect 11056 15258 11080 15260
rect 11136 15258 11160 15260
rect 11216 15258 11240 15260
rect 10976 15206 10986 15258
rect 11230 15206 11240 15258
rect 10976 15204 11000 15206
rect 11056 15204 11080 15206
rect 11136 15204 11160 15206
rect 11216 15204 11240 15206
rect 10920 15195 11296 15204
rect 10920 14172 11296 14181
rect 10976 14170 11000 14172
rect 11056 14170 11080 14172
rect 11136 14170 11160 14172
rect 11216 14170 11240 14172
rect 10976 14118 10986 14170
rect 11230 14118 11240 14170
rect 10976 14116 11000 14118
rect 11056 14116 11080 14118
rect 11136 14116 11160 14118
rect 11216 14116 11240 14118
rect 10920 14107 11296 14116
rect 11348 13326 11376 15864
rect 11624 15722 11652 17274
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11532 15694 11652 15722
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 14618 11468 15438
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 10920 13084 11296 13093
rect 10976 13082 11000 13084
rect 11056 13082 11080 13084
rect 11136 13082 11160 13084
rect 11216 13082 11240 13084
rect 10976 13030 10986 13082
rect 11230 13030 11240 13082
rect 10976 13028 11000 13030
rect 11056 13028 11080 13030
rect 11136 13028 11160 13030
rect 11216 13028 11240 13030
rect 10920 13019 11296 13028
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10704 12838 10824 12866
rect 10704 12442 10732 12838
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10692 12436 10744 12442
rect 10888 12434 10916 12922
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10692 12378 10744 12384
rect 10796 12406 10916 12434
rect 10508 12368 10560 12374
rect 10796 12322 10824 12406
rect 10508 12310 10560 12316
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10428 11558 10456 12106
rect 10520 11898 10548 12310
rect 10612 12294 10824 12322
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10180 11452 10556 11461
rect 10236 11450 10260 11452
rect 10316 11450 10340 11452
rect 10396 11450 10420 11452
rect 10476 11450 10500 11452
rect 10236 11398 10246 11450
rect 10490 11398 10500 11450
rect 10236 11396 10260 11398
rect 10316 11396 10340 11398
rect 10396 11396 10420 11398
rect 10476 11396 10500 11398
rect 10180 11387 10556 11396
rect 10180 10364 10556 10373
rect 10236 10362 10260 10364
rect 10316 10362 10340 10364
rect 10396 10362 10420 10364
rect 10476 10362 10500 10364
rect 10236 10310 10246 10362
rect 10490 10310 10500 10362
rect 10236 10308 10260 10310
rect 10316 10308 10340 10310
rect 10396 10308 10420 10310
rect 10476 10308 10500 10310
rect 10180 10299 10556 10308
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9968 8362 9996 8842
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5914 8984 6258
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5914 9812 6054
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 4180 4924 4556 4933
rect 4236 4922 4260 4924
rect 4316 4922 4340 4924
rect 4396 4922 4420 4924
rect 4476 4922 4500 4924
rect 4236 4870 4246 4922
rect 4490 4870 4500 4922
rect 4236 4868 4260 4870
rect 4316 4868 4340 4870
rect 4396 4868 4420 4870
rect 4476 4868 4500 4870
rect 4180 4859 4556 4868
rect 4920 4380 5296 4389
rect 4976 4378 5000 4380
rect 5056 4378 5080 4380
rect 5136 4378 5160 4380
rect 5216 4378 5240 4380
rect 4976 4326 4986 4378
rect 5230 4326 5240 4378
rect 4976 4324 5000 4326
rect 5056 4324 5080 4326
rect 5136 4324 5160 4326
rect 5216 4324 5240 4326
rect 4920 4315 5296 4324
rect 9232 4146 9260 5170
rect 9324 4826 9352 5170
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9692 4622 9720 5510
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9588 4140 9640 4146
rect 9692 4128 9720 4422
rect 9640 4100 9720 4128
rect 9588 4082 9640 4088
rect 4180 3836 4556 3845
rect 4236 3834 4260 3836
rect 4316 3834 4340 3836
rect 4396 3834 4420 3836
rect 4476 3834 4500 3836
rect 4236 3782 4246 3834
rect 4490 3782 4500 3834
rect 4236 3780 4260 3782
rect 4316 3780 4340 3782
rect 4396 3780 4420 3782
rect 4476 3780 4500 3782
rect 4180 3771 4556 3780
rect 9232 3602 9260 4082
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 9784 3466 9812 4694
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 4920 3292 5296 3301
rect 4976 3290 5000 3292
rect 5056 3290 5080 3292
rect 5136 3290 5160 3292
rect 5216 3290 5240 3292
rect 4976 3238 4986 3290
rect 5230 3238 5240 3290
rect 4976 3236 5000 3238
rect 5056 3236 5080 3238
rect 5136 3236 5160 3238
rect 5216 3236 5240 3238
rect 4920 3227 5296 3236
rect 4180 2748 4556 2757
rect 4236 2746 4260 2748
rect 4316 2746 4340 2748
rect 4396 2746 4420 2748
rect 4476 2746 4500 2748
rect 4236 2694 4246 2746
rect 4490 2694 4500 2746
rect 4236 2692 4260 2694
rect 4316 2692 4340 2694
rect 4396 2692 4420 2694
rect 4476 2692 4500 2694
rect 4180 2683 4556 2692
rect 9876 2650 9904 7822
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9968 6458 9996 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 10060 6322 10088 9454
rect 10180 9276 10556 9285
rect 10236 9274 10260 9276
rect 10316 9274 10340 9276
rect 10396 9274 10420 9276
rect 10476 9274 10500 9276
rect 10236 9222 10246 9274
rect 10490 9222 10500 9274
rect 10236 9220 10260 9222
rect 10316 9220 10340 9222
rect 10396 9220 10420 9222
rect 10476 9220 10500 9222
rect 10180 9211 10556 9220
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8498 10548 8978
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10612 8430 10640 12294
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11354 10732 12174
rect 10784 12096 10836 12102
rect 10980 12084 11008 12854
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10836 12056 11008 12084
rect 11060 12096 11112 12102
rect 10784 12038 10836 12044
rect 11164 12084 11192 12718
rect 11348 12442 11376 13126
rect 11440 12782 11468 14554
rect 11532 13258 11560 15694
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 14482 11652 15574
rect 11716 15026 11744 16526
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12442 11468 12582
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11112 12056 11468 12084
rect 11060 12038 11112 12044
rect 10920 11996 11296 12005
rect 10976 11994 11000 11996
rect 11056 11994 11080 11996
rect 11136 11994 11160 11996
rect 11216 11994 11240 11996
rect 10976 11942 10986 11994
rect 11230 11942 11240 11994
rect 10976 11940 11000 11942
rect 11056 11940 11080 11942
rect 11136 11940 11160 11942
rect 11216 11940 11240 11942
rect 10920 11931 11296 11940
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10704 10674 10732 11290
rect 10888 11218 10916 11834
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11354 11376 11698
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 11440 11082 11468 12056
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 10920 10908 11296 10917
rect 10976 10906 11000 10908
rect 11056 10906 11080 10908
rect 11136 10906 11160 10908
rect 11216 10906 11240 10908
rect 10976 10854 10986 10906
rect 11230 10854 11240 10906
rect 10976 10852 11000 10854
rect 11056 10852 11080 10854
rect 11136 10852 11160 10854
rect 11216 10852 11240 10854
rect 10920 10843 11296 10852
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10920 9820 11296 9829
rect 10976 9818 11000 9820
rect 11056 9818 11080 9820
rect 11136 9818 11160 9820
rect 11216 9818 11240 9820
rect 10976 9766 10986 9818
rect 11230 9766 11240 9818
rect 10976 9764 11000 9766
rect 11056 9764 11080 9766
rect 11136 9764 11160 9766
rect 11216 9764 11240 9766
rect 10920 9755 11296 9764
rect 11532 9602 11560 13194
rect 11624 12918 11652 14418
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11716 12764 11744 14962
rect 11624 12736 11744 12764
rect 11624 12102 11652 12736
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11014 11652 12038
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11164 9574 11560 9602
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9110 11008 9454
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 11072 9042 11100 9522
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11164 8974 11192 9574
rect 11716 9466 11744 12582
rect 11808 12458 11836 21270
rect 11992 20942 12020 21898
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11900 16658 11928 17682
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11900 15434 11928 16390
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14482 11928 14758
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11900 12646 11928 13262
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11808 12430 11928 12458
rect 11900 11626 11928 12430
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 11218 11836 11494
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11348 9438 11744 9466
rect 11348 8974 11376 9438
rect 11520 9376 11572 9382
rect 11808 9364 11836 11018
rect 11520 9318 11572 9324
rect 11716 9336 11836 9364
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 10920 8732 11296 8741
rect 10976 8730 11000 8732
rect 11056 8730 11080 8732
rect 11136 8730 11160 8732
rect 11216 8730 11240 8732
rect 10976 8678 10986 8730
rect 11230 8678 11240 8730
rect 10976 8676 11000 8678
rect 11056 8676 11080 8678
rect 11136 8676 11160 8678
rect 11216 8676 11240 8678
rect 10920 8667 11296 8676
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 11348 8378 11376 8910
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11440 8480 11468 8774
rect 11532 8634 11560 9318
rect 11716 8838 11744 9336
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11440 8452 11560 8480
rect 10180 8188 10556 8197
rect 10236 8186 10260 8188
rect 10316 8186 10340 8188
rect 10396 8186 10420 8188
rect 10476 8186 10500 8188
rect 10236 8134 10246 8186
rect 10490 8134 10500 8186
rect 10236 8132 10260 8134
rect 10316 8132 10340 8134
rect 10396 8132 10420 8134
rect 10476 8132 10500 8134
rect 10180 8123 10556 8132
rect 10180 7100 10556 7109
rect 10236 7098 10260 7100
rect 10316 7098 10340 7100
rect 10396 7098 10420 7100
rect 10476 7098 10500 7100
rect 10236 7046 10246 7098
rect 10490 7046 10500 7098
rect 10236 7044 10260 7046
rect 10316 7044 10340 7046
rect 10396 7044 10420 7046
rect 10476 7044 10500 7046
rect 10180 7035 10556 7044
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10612 6202 10640 8366
rect 11348 8350 11468 8378
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 7886 11376 8230
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 10920 7644 11296 7653
rect 10976 7642 11000 7644
rect 11056 7642 11080 7644
rect 11136 7642 11160 7644
rect 11216 7642 11240 7644
rect 10976 7590 10986 7642
rect 11230 7590 11240 7642
rect 10976 7588 11000 7590
rect 11056 7588 11080 7590
rect 11136 7588 11160 7590
rect 11216 7588 11240 7590
rect 10920 7579 11296 7588
rect 11440 6798 11468 8350
rect 11532 6798 11560 8452
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6254 10824 6666
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 10920 6556 11296 6565
rect 10976 6554 11000 6556
rect 11056 6554 11080 6556
rect 11136 6554 11160 6556
rect 11216 6554 11240 6556
rect 10976 6502 10986 6554
rect 11230 6502 11240 6554
rect 10976 6500 11000 6502
rect 11056 6500 11080 6502
rect 11136 6500 11160 6502
rect 11216 6500 11240 6502
rect 10920 6491 11296 6500
rect 10784 6248 10836 6254
rect 10612 6174 10732 6202
rect 10784 6190 10836 6196
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10180 6012 10556 6021
rect 10236 6010 10260 6012
rect 10316 6010 10340 6012
rect 10396 6010 10420 6012
rect 10476 6010 10500 6012
rect 10236 5958 10246 6010
rect 10490 5958 10500 6010
rect 10236 5956 10260 5958
rect 10316 5956 10340 5958
rect 10396 5956 10420 5958
rect 10476 5956 10500 5958
rect 10180 5947 10556 5956
rect 10612 5914 10640 6054
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10704 5778 10732 6174
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5012 10180 5510
rect 10060 4984 10180 5012
rect 10060 4622 10088 4984
rect 10180 4924 10556 4933
rect 10236 4922 10260 4924
rect 10316 4922 10340 4924
rect 10396 4922 10420 4924
rect 10476 4922 10500 4924
rect 10236 4870 10246 4922
rect 10490 4870 10500 4922
rect 10236 4868 10260 4870
rect 10316 4868 10340 4870
rect 10396 4868 10420 4870
rect 10476 4868 10500 4870
rect 10180 4859 10556 4868
rect 10612 4622 10640 5578
rect 10796 5370 10824 6190
rect 11348 5710 11376 6598
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11624 5914 11652 6190
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5794 11744 8774
rect 11808 8634 11836 8774
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11992 6322 12020 19654
rect 12084 12238 12112 22066
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12544 21146 12572 21490
rect 12532 21140 12584 21146
rect 12532 21082 12584 21088
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12268 20482 12296 20742
rect 12636 20602 12664 20878
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12176 20466 12296 20482
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12164 20460 12296 20466
rect 12216 20454 12296 20460
rect 12164 20402 12216 20408
rect 12452 18290 12480 20470
rect 12728 20058 12756 22066
rect 13268 22034 13320 22040
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21690 13124 21966
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 13004 21078 13032 21422
rect 13096 21146 13124 21626
rect 13176 21344 13228 21350
rect 13176 21286 13228 21292
rect 13188 21146 13216 21286
rect 13280 21146 13308 22034
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 13648 20398 13676 21422
rect 13740 21010 13768 22510
rect 14096 22160 14148 22166
rect 14096 22102 14148 22108
rect 14108 21690 14136 22102
rect 14476 21962 14504 22578
rect 14464 21956 14516 21962
rect 14464 21898 14516 21904
rect 14096 21684 14148 21690
rect 14096 21626 14148 21632
rect 14568 21486 14596 23598
rect 14752 22710 14780 25638
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14936 24410 14964 24686
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14936 22778 14964 24346
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15120 23866 15148 24142
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14752 21350 14780 22646
rect 15120 22642 15148 23802
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15212 22574 15240 26454
rect 15304 26450 15332 29242
rect 15396 28558 15424 29514
rect 16040 29510 16068 29582
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 16132 29306 16160 29446
rect 16920 29404 17296 29413
rect 16976 29402 17000 29404
rect 17056 29402 17080 29404
rect 17136 29402 17160 29404
rect 17216 29402 17240 29404
rect 16976 29350 16986 29402
rect 17230 29350 17240 29402
rect 16976 29348 17000 29350
rect 17056 29348 17080 29350
rect 17136 29348 17160 29350
rect 17216 29348 17240 29350
rect 16920 29339 17296 29348
rect 16120 29300 16172 29306
rect 16120 29242 16172 29248
rect 16180 28860 16556 28869
rect 16236 28858 16260 28860
rect 16316 28858 16340 28860
rect 16396 28858 16420 28860
rect 16476 28858 16500 28860
rect 16236 28806 16246 28858
rect 16490 28806 16500 28858
rect 16236 28804 16260 28806
rect 16316 28804 16340 28806
rect 16396 28804 16420 28806
rect 16476 28804 16500 28806
rect 16180 28795 16556 28804
rect 17328 28558 17356 29582
rect 17972 29050 18000 29990
rect 17880 29022 18000 29050
rect 17684 28960 17736 28966
rect 17684 28902 17736 28908
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 15568 28484 15620 28490
rect 15568 28426 15620 28432
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15212 21622 15240 22170
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13740 20466 13768 20946
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14108 20602 14136 20742
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14660 20466 14688 20878
rect 14752 20466 14780 21286
rect 15304 20874 15332 24006
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12728 19922 12756 19994
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 14016 19854 14044 20266
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14200 19514 14228 20334
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14844 19446 14872 20402
rect 15304 19922 15332 20810
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 14832 19440 14884 19446
rect 14832 19382 14884 19388
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15108 18896 15160 18902
rect 15108 18838 15160 18844
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14188 18760 14240 18766
rect 14740 18760 14792 18766
rect 14188 18702 14240 18708
rect 14738 18728 14740 18737
rect 14792 18728 14794 18737
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18358 12756 18566
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12268 17785 12296 17818
rect 12254 17776 12310 17785
rect 12452 17746 12480 18226
rect 14108 17882 14136 18702
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 12254 17711 12310 17720
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17338 12204 17614
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 13648 17134 13676 17682
rect 14096 17604 14148 17610
rect 14096 17546 14148 17552
rect 13452 17128 13504 17134
rect 13450 17096 13452 17105
rect 13636 17128 13688 17134
rect 13504 17096 13506 17105
rect 13636 17070 13688 17076
rect 13450 17031 13506 17040
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15502 12204 15846
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14006 12204 14758
rect 12268 14006 12296 16934
rect 14108 16794 14136 17546
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14200 16522 14228 18702
rect 14738 18663 14794 18672
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14292 16674 14320 18158
rect 15120 18086 15148 18838
rect 15212 18290 15240 19178
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 14568 17746 14596 18022
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14384 17202 14412 17478
rect 14476 17377 14504 17478
rect 14462 17368 14518 17377
rect 14462 17303 14518 17312
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14384 16794 14412 17138
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14292 16646 14412 16674
rect 14384 16522 14412 16646
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12636 15162 12664 16050
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14074 12480 14894
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12256 12232 12308 12238
rect 12360 12186 12388 13942
rect 12820 13938 12848 15846
rect 13280 15706 13308 15982
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13188 15162 13216 15642
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15162 14136 15302
rect 14476 15162 14504 17303
rect 14752 17241 14780 17682
rect 15120 17270 15148 18022
rect 15200 17808 15252 17814
rect 15198 17776 15200 17785
rect 15252 17776 15254 17785
rect 15198 17711 15254 17720
rect 15198 17368 15254 17377
rect 15198 17303 15200 17312
rect 15252 17303 15254 17312
rect 15200 17274 15252 17280
rect 15108 17264 15160 17270
rect 14738 17232 14794 17241
rect 15108 17206 15160 17212
rect 14738 17167 14794 17176
rect 15304 16658 15332 19450
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 15978 14780 16526
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13464 14482 13492 14894
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12308 12180 12388 12186
rect 12256 12174 12388 12180
rect 12268 12158 12388 12174
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11898 12112 12038
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 8974 12112 10950
rect 12176 9586 12204 11086
rect 12268 9586 12296 11562
rect 12360 9602 12388 12158
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11218 12572 11494
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12728 11082 12756 12038
rect 12912 11626 12940 13330
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12256 9580 12308 9586
rect 12360 9574 12480 9602
rect 12256 9522 12308 9528
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11624 5766 11744 5794
rect 11624 5710 11652 5766
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 10920 5468 11296 5477
rect 10976 5466 11000 5468
rect 11056 5466 11080 5468
rect 11136 5466 11160 5468
rect 11216 5466 11240 5468
rect 10976 5414 10986 5466
rect 11230 5414 11240 5466
rect 10976 5412 11000 5414
rect 11056 5412 11080 5414
rect 11136 5412 11160 5414
rect 11216 5412 11240 5414
rect 10920 5403 11296 5412
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 11440 5166 11468 5646
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11532 5370 11560 5510
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10180 3836 10556 3845
rect 10236 3834 10260 3836
rect 10316 3834 10340 3836
rect 10396 3834 10420 3836
rect 10476 3834 10500 3836
rect 10236 3782 10246 3834
rect 10490 3782 10500 3834
rect 10236 3780 10260 3782
rect 10316 3780 10340 3782
rect 10396 3780 10420 3782
rect 10476 3780 10500 3782
rect 10180 3771 10556 3780
rect 10704 3738 10732 4422
rect 10920 4380 11296 4389
rect 10976 4378 11000 4380
rect 11056 4378 11080 4380
rect 11136 4378 11160 4380
rect 11216 4378 11240 4380
rect 10976 4326 10986 4378
rect 11230 4326 11240 4378
rect 10976 4324 11000 4326
rect 11056 4324 11080 4326
rect 11136 4324 11160 4326
rect 11216 4324 11240 4326
rect 10920 4315 11296 4324
rect 11440 4010 11468 5102
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 11716 3602 11744 5578
rect 11900 4622 11928 6054
rect 12084 5710 12112 8910
rect 12176 8634 12204 9522
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9178 12388 9454
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12452 9058 12480 9574
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12360 9030 12480 9058
rect 12532 9036 12584 9042
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12176 7886 12204 8570
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12360 5302 12388 9030
rect 12532 8978 12584 8984
rect 12544 8498 12572 8978
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 5370 12664 9318
rect 12912 9042 12940 11562
rect 13188 11558 13216 12718
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12084 4622 12112 5238
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12452 4146 12480 4966
rect 12636 4826 12664 5170
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 11900 3738 11928 4082
rect 12544 3738 12572 4490
rect 12912 4486 12940 8978
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 13004 3602 13032 4422
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 10920 3292 11296 3301
rect 10976 3290 11000 3292
rect 11056 3290 11080 3292
rect 11136 3290 11160 3292
rect 11216 3290 11240 3292
rect 10976 3238 10986 3290
rect 11230 3238 11240 3290
rect 10976 3236 11000 3238
rect 11056 3236 11080 3238
rect 11136 3236 11160 3238
rect 11216 3236 11240 3238
rect 10920 3227 11296 3236
rect 10180 2748 10556 2757
rect 10236 2746 10260 2748
rect 10316 2746 10340 2748
rect 10396 2746 10420 2748
rect 10476 2746 10500 2748
rect 10236 2694 10246 2746
rect 10490 2694 10500 2746
rect 10236 2692 10260 2694
rect 10316 2692 10340 2694
rect 10396 2692 10420 2694
rect 10476 2692 10500 2694
rect 10180 2683 10556 2692
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10796 2378 10916 2394
rect 13280 2378 13308 14214
rect 13464 12434 13492 14418
rect 13648 14278 13676 14894
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14414 13768 14758
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13924 14346 13952 14486
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14108 13530 14136 13874
rect 14200 13870 14228 14350
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14096 12912 14148 12918
rect 14200 12900 14228 13806
rect 14476 13326 14504 15098
rect 14752 14958 14780 15914
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 14740 14952 14792 14958
rect 14660 14912 14740 14940
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14660 13258 14688 14912
rect 14740 14894 14792 14900
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14148 12872 14228 12900
rect 14096 12854 14148 12860
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13464 12406 13676 12434
rect 13464 12374 13492 12406
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13372 8634 13400 8842
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13556 5778 13584 8366
rect 13648 6236 13676 12406
rect 13740 12306 13768 12582
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13832 11898 13860 12038
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14108 11762 14136 12854
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 11898 14228 12106
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14096 11620 14148 11626
rect 14280 11620 14332 11626
rect 14148 11580 14280 11608
rect 14096 11562 14148 11568
rect 14280 11562 14332 11568
rect 14660 9674 14688 13194
rect 14844 11762 14872 15846
rect 15120 15706 15148 15846
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 15212 15026 15240 16390
rect 15396 15638 15424 28358
rect 15580 28218 15608 28426
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 15764 27674 15792 28494
rect 16920 28316 17296 28325
rect 16976 28314 17000 28316
rect 17056 28314 17080 28316
rect 17136 28314 17160 28316
rect 17216 28314 17240 28316
rect 16976 28262 16986 28314
rect 17230 28262 17240 28314
rect 16976 28260 17000 28262
rect 17056 28260 17080 28262
rect 17136 28260 17160 28262
rect 17216 28260 17240 28262
rect 16920 28251 17296 28260
rect 17328 28014 17356 28494
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 17512 28218 17540 28426
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17696 28150 17724 28902
rect 17684 28144 17736 28150
rect 17684 28086 17736 28092
rect 17316 28008 17368 28014
rect 17316 27950 17368 27956
rect 16180 27772 16556 27781
rect 16236 27770 16260 27772
rect 16316 27770 16340 27772
rect 16396 27770 16420 27772
rect 16476 27770 16500 27772
rect 16236 27718 16246 27770
rect 16490 27718 16500 27770
rect 16236 27716 16260 27718
rect 16316 27716 16340 27718
rect 16396 27716 16420 27718
rect 16476 27716 16500 27718
rect 16180 27707 16556 27716
rect 15752 27668 15804 27674
rect 15752 27610 15804 27616
rect 16580 27600 16632 27606
rect 16580 27542 16632 27548
rect 16592 27470 16620 27542
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 16580 27464 16632 27470
rect 16580 27406 16632 27412
rect 15764 27130 15792 27406
rect 16672 27396 16724 27402
rect 16672 27338 16724 27344
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 16040 26450 16068 27270
rect 16180 26684 16556 26693
rect 16236 26682 16260 26684
rect 16316 26682 16340 26684
rect 16396 26682 16420 26684
rect 16476 26682 16500 26684
rect 16236 26630 16246 26682
rect 16490 26630 16500 26682
rect 16236 26628 16260 26630
rect 16316 26628 16340 26630
rect 16396 26628 16420 26630
rect 16476 26628 16500 26630
rect 16180 26619 16556 26628
rect 16684 26586 16712 27338
rect 16856 27328 16908 27334
rect 16776 27288 16856 27316
rect 16776 27062 16804 27288
rect 16856 27270 16908 27276
rect 16920 27228 17296 27237
rect 16976 27226 17000 27228
rect 17056 27226 17080 27228
rect 17136 27226 17160 27228
rect 17216 27226 17240 27228
rect 16976 27174 16986 27226
rect 17230 27174 17240 27226
rect 16976 27172 17000 27174
rect 17056 27172 17080 27174
rect 17136 27172 17160 27174
rect 17216 27172 17240 27174
rect 16920 27163 17296 27172
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 17328 26926 17356 27950
rect 17040 26920 17092 26926
rect 17040 26862 17092 26868
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 17052 26450 17080 26862
rect 16028 26444 16080 26450
rect 16028 26386 16080 26392
rect 17040 26444 17092 26450
rect 17040 26386 17092 26392
rect 16920 26140 17296 26149
rect 16976 26138 17000 26140
rect 17056 26138 17080 26140
rect 17136 26138 17160 26140
rect 17216 26138 17240 26140
rect 16976 26086 16986 26138
rect 17230 26086 17240 26138
rect 16976 26084 17000 26086
rect 17056 26084 17080 26086
rect 17136 26084 17160 26086
rect 17216 26084 17240 26086
rect 16920 26075 17296 26084
rect 16180 25596 16556 25605
rect 16236 25594 16260 25596
rect 16316 25594 16340 25596
rect 16396 25594 16420 25596
rect 16476 25594 16500 25596
rect 16236 25542 16246 25594
rect 16490 25542 16500 25594
rect 16236 25540 16260 25542
rect 16316 25540 16340 25542
rect 16396 25540 16420 25542
rect 16476 25540 16500 25542
rect 16180 25531 16556 25540
rect 17880 25362 17908 29022
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17972 25906 18000 26182
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 16920 25052 17296 25061
rect 16976 25050 17000 25052
rect 17056 25050 17080 25052
rect 17136 25050 17160 25052
rect 17216 25050 17240 25052
rect 16976 24998 16986 25050
rect 17230 24998 17240 25050
rect 16976 24996 17000 24998
rect 17056 24996 17080 24998
rect 17136 24996 17160 24998
rect 17216 24996 17240 24998
rect 16920 24987 17296 24996
rect 17512 24954 17540 25094
rect 17500 24948 17552 24954
rect 17880 24936 17908 25298
rect 17500 24890 17552 24896
rect 17788 24908 17908 24936
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17224 24608 17276 24614
rect 17224 24550 17276 24556
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 16180 24508 16556 24517
rect 16236 24506 16260 24508
rect 16316 24506 16340 24508
rect 16396 24506 16420 24508
rect 16476 24506 16500 24508
rect 16236 24454 16246 24506
rect 16490 24454 16500 24506
rect 16236 24452 16260 24454
rect 16316 24452 16340 24454
rect 16396 24452 16420 24454
rect 16476 24452 16500 24454
rect 16180 24443 16556 24452
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 15488 22234 15516 23122
rect 15764 23118 15792 24006
rect 16132 23866 16160 24210
rect 17236 24138 17264 24550
rect 17512 24138 17540 24550
rect 17224 24132 17276 24138
rect 17224 24074 17276 24080
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 16920 23964 17296 23973
rect 16976 23962 17000 23964
rect 17056 23962 17080 23964
rect 17136 23962 17160 23964
rect 17216 23962 17240 23964
rect 16976 23910 16986 23962
rect 17230 23910 17240 23962
rect 16976 23908 17000 23910
rect 17056 23908 17080 23910
rect 17136 23908 17160 23910
rect 17216 23908 17240 23910
rect 16920 23899 17296 23908
rect 17604 23866 17632 24754
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 16224 23508 16252 23666
rect 17236 23633 17264 23666
rect 17222 23624 17278 23633
rect 17222 23559 17278 23568
rect 16040 23480 16252 23508
rect 16040 23322 16068 23480
rect 16180 23420 16556 23429
rect 16236 23418 16260 23420
rect 16316 23418 16340 23420
rect 16396 23418 16420 23420
rect 16476 23418 16500 23420
rect 16236 23366 16246 23418
rect 16490 23366 16500 23418
rect 16236 23364 16260 23366
rect 16316 23364 16340 23366
rect 16396 23364 16420 23366
rect 16476 23364 16500 23366
rect 16180 23355 16556 23364
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 17788 23186 17816 24908
rect 17972 24834 18000 25842
rect 17880 24806 18000 24834
rect 17880 23798 17908 24806
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17880 23497 17908 23734
rect 17866 23488 17922 23497
rect 17866 23423 17922 23432
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 16920 22876 17296 22885
rect 16976 22874 17000 22876
rect 17056 22874 17080 22876
rect 17136 22874 17160 22876
rect 17216 22874 17240 22876
rect 16976 22822 16986 22874
rect 17230 22822 17240 22874
rect 16976 22820 17000 22822
rect 17056 22820 17080 22822
rect 17136 22820 17160 22822
rect 17216 22820 17240 22822
rect 16920 22811 17296 22820
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16180 22332 16556 22341
rect 16236 22330 16260 22332
rect 16316 22330 16340 22332
rect 16396 22330 16420 22332
rect 16476 22330 16500 22332
rect 16236 22278 16246 22330
rect 16490 22278 16500 22330
rect 16236 22276 16260 22278
rect 16316 22276 16340 22278
rect 16396 22276 16420 22278
rect 16476 22276 16500 22278
rect 16180 22267 16556 22276
rect 15476 22228 15528 22234
rect 15476 22170 15528 22176
rect 16580 22160 16632 22166
rect 16580 22102 16632 22108
rect 16486 21992 16542 22001
rect 16120 21956 16172 21962
rect 16040 21916 16120 21944
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 21690 15884 21830
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 21078 15884 21422
rect 15844 21072 15896 21078
rect 15844 21014 15896 21020
rect 16040 21026 16068 21916
rect 16120 21898 16172 21904
rect 16304 21956 16356 21962
rect 16486 21927 16488 21936
rect 16304 21898 16356 21904
rect 16540 21927 16542 21936
rect 16488 21898 16540 21904
rect 16316 21554 16344 21898
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16488 21480 16540 21486
rect 16592 21468 16620 22102
rect 16540 21440 16620 21468
rect 16488 21422 16540 21428
rect 16500 21350 16528 21422
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16180 21244 16556 21253
rect 16236 21242 16260 21244
rect 16316 21242 16340 21244
rect 16396 21242 16420 21244
rect 16476 21242 16500 21244
rect 16236 21190 16246 21242
rect 16490 21190 16500 21242
rect 16236 21188 16260 21190
rect 16316 21188 16340 21190
rect 16396 21188 16420 21190
rect 16476 21188 16500 21190
rect 16180 21179 16556 21188
rect 16040 20998 16160 21026
rect 16776 21010 16804 22442
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16960 22030 16988 22374
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17406 21992 17462 22001
rect 17406 21927 17462 21936
rect 16920 21788 17296 21797
rect 16976 21786 17000 21788
rect 17056 21786 17080 21788
rect 17136 21786 17160 21788
rect 17216 21786 17240 21788
rect 16976 21734 16986 21786
rect 17230 21734 17240 21786
rect 16976 21732 17000 21734
rect 17056 21732 17080 21734
rect 17136 21732 17160 21734
rect 17216 21732 17240 21734
rect 16920 21723 17296 21732
rect 17420 21690 17448 21927
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16960 21010 16988 21558
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16040 20602 16068 20878
rect 16132 20602 16160 20998
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15474 19408 15530 19417
rect 15580 19378 15608 20402
rect 16040 20346 16068 20402
rect 16500 20398 16528 20878
rect 16684 20534 16712 20946
rect 16960 20913 16988 20946
rect 16946 20904 17002 20913
rect 16946 20839 17002 20848
rect 17144 20806 17172 21490
rect 17224 21480 17276 21486
rect 17224 21422 17276 21428
rect 17236 21146 17264 21422
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 16920 20700 17296 20709
rect 16976 20698 17000 20700
rect 17056 20698 17080 20700
rect 17136 20698 17160 20700
rect 17216 20698 17240 20700
rect 16976 20646 16986 20698
rect 17230 20646 17240 20698
rect 16976 20644 17000 20646
rect 17056 20644 17080 20646
rect 17136 20644 17160 20646
rect 17216 20644 17240 20646
rect 16920 20635 17296 20644
rect 16672 20528 16724 20534
rect 16724 20488 16804 20516
rect 16672 20470 16724 20476
rect 15948 20318 16068 20346
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15764 19446 15792 19926
rect 15856 19446 15884 20198
rect 15948 19961 15976 20318
rect 16028 20256 16080 20262
rect 16500 20244 16528 20334
rect 16500 20216 16620 20244
rect 16028 20198 16080 20204
rect 15934 19952 15990 19961
rect 15934 19887 15990 19896
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15752 19440 15804 19446
rect 15752 19382 15804 19388
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15474 19343 15530 19352
rect 15568 19372 15620 19378
rect 15488 19174 15516 19343
rect 15568 19314 15620 19320
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15488 17746 15516 18158
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15304 15162 15332 15302
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15304 14618 15332 14826
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14752 11354 14780 11698
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14384 9646 14688 9674
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8498 13860 8978
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13832 6458 13860 8434
rect 14384 8430 14412 9646
rect 14844 9058 14872 11698
rect 15120 11150 15148 13874
rect 15488 13530 15516 17682
rect 15580 17610 15608 19314
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 18834 15700 19110
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15764 18442 15792 19382
rect 15764 18414 15884 18442
rect 15948 18426 15976 19790
rect 16040 19718 16068 20198
rect 16180 20156 16556 20165
rect 16236 20154 16260 20156
rect 16316 20154 16340 20156
rect 16396 20154 16420 20156
rect 16476 20154 16500 20156
rect 16236 20102 16246 20154
rect 16490 20102 16500 20154
rect 16236 20100 16260 20102
rect 16316 20100 16340 20102
rect 16396 20100 16420 20102
rect 16476 20100 16500 20102
rect 16180 20091 16556 20100
rect 16592 20040 16620 20216
rect 16500 20012 16620 20040
rect 16672 20052 16724 20058
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 16500 19514 16528 20012
rect 16672 19994 16724 20000
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16180 19068 16556 19077
rect 16236 19066 16260 19068
rect 16316 19066 16340 19068
rect 16396 19066 16420 19068
rect 16476 19066 16500 19068
rect 16236 19014 16246 19066
rect 16490 19014 16500 19066
rect 16236 19012 16260 19014
rect 16316 19012 16340 19014
rect 16396 19012 16420 19014
rect 16476 19012 16500 19014
rect 16180 19003 16556 19012
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16316 18873 16344 18906
rect 16302 18864 16358 18873
rect 16302 18799 16358 18808
rect 16488 18828 16540 18834
rect 15856 18358 15884 18414
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 18352 15896 18358
rect 15844 18294 15896 18300
rect 16316 18290 16344 18799
rect 16488 18770 16540 18776
rect 16500 18358 16528 18770
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15948 17814 15976 18158
rect 15936 17808 15988 17814
rect 15934 17776 15936 17785
rect 15988 17776 15990 17785
rect 15660 17740 15712 17746
rect 15934 17711 15990 17720
rect 15660 17682 15712 17688
rect 15672 17649 15700 17682
rect 15658 17640 15714 17649
rect 15568 17604 15620 17610
rect 15658 17575 15714 17584
rect 15752 17604 15804 17610
rect 15568 17546 15620 17552
rect 15752 17546 15804 17552
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16250 15700 16458
rect 15764 16454 15792 17546
rect 15948 16794 15976 17546
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16040 16590 16068 18226
rect 16592 18222 16620 19246
rect 16684 18426 16712 19994
rect 16776 19854 16804 20488
rect 17512 20262 17540 20946
rect 17604 20534 17632 22102
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17696 20806 17724 20878
rect 17684 20800 17736 20806
rect 17684 20742 17736 20748
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 16920 19612 17296 19621
rect 16976 19610 17000 19612
rect 17056 19610 17080 19612
rect 17136 19610 17160 19612
rect 17216 19610 17240 19612
rect 16976 19558 16986 19610
rect 17230 19558 17240 19610
rect 16976 19556 17000 19558
rect 17056 19556 17080 19558
rect 17136 19556 17160 19558
rect 17216 19556 17240 19558
rect 16920 19547 17296 19556
rect 16946 19408 17002 19417
rect 17420 19378 17448 19790
rect 17512 19786 17540 20198
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 16946 19343 17002 19352
rect 17408 19372 17460 19378
rect 16960 18834 16988 19343
rect 17408 19314 17460 19320
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 18442 16804 18702
rect 16920 18524 17296 18533
rect 16976 18522 17000 18524
rect 17056 18522 17080 18524
rect 17136 18522 17160 18524
rect 17216 18522 17240 18524
rect 16976 18470 16986 18522
rect 17230 18470 17240 18522
rect 16976 18468 17000 18470
rect 17056 18468 17080 18470
rect 17136 18468 17160 18470
rect 17216 18468 17240 18470
rect 16920 18459 17296 18468
rect 16672 18420 16724 18426
rect 16776 18414 16896 18442
rect 16672 18362 16724 18368
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16180 17980 16556 17989
rect 16236 17978 16260 17980
rect 16316 17978 16340 17980
rect 16396 17978 16420 17980
rect 16476 17978 16500 17980
rect 16236 17926 16246 17978
rect 16490 17926 16500 17978
rect 16236 17924 16260 17926
rect 16316 17924 16340 17926
rect 16396 17924 16420 17926
rect 16476 17924 16500 17926
rect 16180 17915 16556 17924
rect 16486 17232 16542 17241
rect 16486 17167 16488 17176
rect 16540 17167 16542 17176
rect 16488 17138 16540 17144
rect 16592 17134 16620 18158
rect 16684 17338 16712 18362
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16776 17746 16804 18294
rect 16868 18290 16896 18414
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 16868 17814 16896 18226
rect 17236 17882 17264 18226
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 17328 17649 17356 19178
rect 17420 18834 17448 19314
rect 17512 18834 17540 19722
rect 17696 19378 17724 20742
rect 17788 20466 17816 21422
rect 17880 21146 17908 21490
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17880 20466 17908 21082
rect 18064 20942 18092 21558
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18064 20602 18092 20878
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17788 20262 17816 20402
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17408 18692 17460 18698
rect 17408 18634 17460 18640
rect 17314 17640 17370 17649
rect 17314 17575 17370 17584
rect 16920 17436 17296 17445
rect 16976 17434 17000 17436
rect 17056 17434 17080 17436
rect 17136 17434 17160 17436
rect 17216 17434 17240 17436
rect 16976 17382 16986 17434
rect 17230 17382 17240 17434
rect 16976 17380 17000 17382
rect 17056 17380 17080 17382
rect 17136 17380 17160 17382
rect 17216 17380 17240 17382
rect 16920 17371 17296 17380
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16776 16998 16804 17206
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16180 16892 16556 16901
rect 16236 16890 16260 16892
rect 16316 16890 16340 16892
rect 16396 16890 16420 16892
rect 16476 16890 16500 16892
rect 16236 16838 16246 16890
rect 16490 16838 16500 16890
rect 16236 16836 16260 16838
rect 16316 16836 16340 16838
rect 16396 16836 16420 16838
rect 16476 16836 16500 16838
rect 16180 16827 16556 16836
rect 16684 16794 16712 16934
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 16776 16250 16804 16934
rect 16920 16348 17296 16357
rect 16976 16346 17000 16348
rect 17056 16346 17080 16348
rect 17136 16346 17160 16348
rect 17216 16346 17240 16348
rect 16976 16294 16986 16346
rect 17230 16294 17240 16346
rect 16976 16292 17000 16294
rect 17056 16292 17080 16294
rect 17136 16292 17160 16294
rect 17216 16292 17240 16294
rect 16920 16283 17296 16292
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15580 15026 15608 15438
rect 15672 15026 15700 16186
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15580 14618 15608 14962
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15764 14074 15792 14962
rect 15948 14906 15976 15098
rect 15856 14878 15976 14906
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15764 13938 15792 14010
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15856 13818 15884 14878
rect 15764 13790 15884 13818
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15212 13190 15240 13262
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15396 11898 15424 12174
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14844 9030 14964 9058
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14844 7886 14872 8842
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7546 14688 7686
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14844 7410 14872 7822
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13820 6248 13872 6254
rect 13648 6208 13820 6236
rect 13820 6190 13872 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5914 13676 6054
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4758 13860 4966
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13924 4162 13952 5102
rect 14200 5030 14228 6122
rect 14844 5710 14872 7346
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14108 4826 14136 4966
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14200 4622 14228 4966
rect 14384 4622 14412 5102
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 13832 4146 13952 4162
rect 13820 4140 13952 4146
rect 13872 4134 13952 4140
rect 13820 4082 13872 4088
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13372 2514 13400 4014
rect 14384 3942 14412 4558
rect 14844 4078 14872 5646
rect 14936 5098 14964 9030
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 15028 7886 15056 8230
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15200 6248 15252 6254
rect 15200 6190 15252 6196
rect 15212 5914 15240 6190
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15212 5234 15240 5850
rect 15304 5370 15332 11630
rect 15382 11112 15438 11121
rect 15382 11047 15438 11056
rect 15396 9654 15424 11047
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 8634 15516 8774
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14936 4826 14964 5034
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 15304 4622 15332 5306
rect 15764 4706 15792 13790
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13394 15884 13670
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15856 4842 15884 13126
rect 16040 11762 16068 16118
rect 16180 15804 16556 15813
rect 16236 15802 16260 15804
rect 16316 15802 16340 15804
rect 16396 15802 16420 15804
rect 16476 15802 16500 15804
rect 16236 15750 16246 15802
rect 16490 15750 16500 15802
rect 16236 15748 16260 15750
rect 16316 15748 16340 15750
rect 16396 15748 16420 15750
rect 16476 15748 16500 15750
rect 16180 15739 16556 15748
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 16132 15026 16160 15574
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15094 16252 15302
rect 16920 15260 17296 15269
rect 16976 15258 17000 15260
rect 17056 15258 17080 15260
rect 17136 15258 17160 15260
rect 17216 15258 17240 15260
rect 16976 15206 16986 15258
rect 17230 15206 17240 15258
rect 16976 15204 17000 15206
rect 17056 15204 17080 15206
rect 17136 15204 17160 15206
rect 17216 15204 17240 15206
rect 16920 15195 17296 15204
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16180 14716 16556 14725
rect 16236 14714 16260 14716
rect 16316 14714 16340 14716
rect 16396 14714 16420 14716
rect 16476 14714 16500 14716
rect 16236 14662 16246 14714
rect 16490 14662 16500 14714
rect 16236 14660 16260 14662
rect 16316 14660 16340 14662
rect 16396 14660 16420 14662
rect 16476 14660 16500 14662
rect 16180 14651 16556 14660
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 14226 16896 14350
rect 16776 14198 16896 14226
rect 16180 13628 16556 13637
rect 16236 13626 16260 13628
rect 16316 13626 16340 13628
rect 16396 13626 16420 13628
rect 16476 13626 16500 13628
rect 16236 13574 16246 13626
rect 16490 13574 16500 13626
rect 16236 13572 16260 13574
rect 16316 13572 16340 13574
rect 16396 13572 16420 13574
rect 16476 13572 16500 13574
rect 16180 13563 16556 13572
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16132 13326 16160 13466
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16180 12540 16556 12549
rect 16236 12538 16260 12540
rect 16316 12538 16340 12540
rect 16396 12538 16420 12540
rect 16476 12538 16500 12540
rect 16236 12486 16246 12538
rect 16490 12486 16500 12538
rect 16236 12484 16260 12486
rect 16316 12484 16340 12486
rect 16396 12484 16420 12486
rect 16476 12484 16500 12486
rect 16180 12475 16556 12484
rect 16684 12434 16712 12582
rect 16592 12406 16712 12434
rect 16592 11762 16620 12406
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11898 16712 12038
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16776 11830 16804 14198
rect 16920 14172 17296 14181
rect 16976 14170 17000 14172
rect 17056 14170 17080 14172
rect 17136 14170 17160 14172
rect 17216 14170 17240 14172
rect 16976 14118 16986 14170
rect 17230 14118 17240 14170
rect 16976 14116 17000 14118
rect 17056 14116 17080 14118
rect 17136 14116 17160 14118
rect 17216 14116 17240 14118
rect 16920 14107 17296 14116
rect 16920 13084 17296 13093
rect 16976 13082 17000 13084
rect 17056 13082 17080 13084
rect 17136 13082 17160 13084
rect 17216 13082 17240 13084
rect 16976 13030 16986 13082
rect 17230 13030 17240 13082
rect 16976 13028 17000 13030
rect 17056 13028 17080 13030
rect 17136 13028 17160 13030
rect 17216 13028 17240 13030
rect 16920 13019 17296 13028
rect 17328 12986 17356 17575
rect 17420 17066 17448 18634
rect 17512 18222 17540 18770
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 17746 17540 18158
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17604 17082 17632 19110
rect 17696 18630 17724 19314
rect 17880 18766 17908 20198
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17868 18760 17920 18766
rect 17972 18737 18000 18770
rect 17868 18702 17920 18708
rect 17958 18728 18014 18737
rect 17958 18663 18014 18672
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 17270 17724 18566
rect 17776 18216 17828 18222
rect 17776 18158 17828 18164
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17408 17060 17460 17066
rect 17604 17054 17724 17082
rect 17408 17002 17460 17008
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12442 17080 12786
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17144 12102 17172 12718
rect 17420 12434 17448 17002
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 14482 17540 14758
rect 17604 14618 17632 16662
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17328 12406 17448 12434
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 16920 11996 17296 12005
rect 16976 11994 17000 11996
rect 17056 11994 17080 11996
rect 17136 11994 17160 11996
rect 17216 11994 17240 11996
rect 16976 11942 16986 11994
rect 17230 11942 17240 11994
rect 16976 11940 17000 11942
rect 17056 11940 17080 11942
rect 17136 11940 17160 11942
rect 17216 11940 17240 11942
rect 16920 11931 17296 11940
rect 17328 11880 17356 12406
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17236 11852 17356 11880
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11082 16068 11494
rect 16180 11452 16556 11461
rect 16236 11450 16260 11452
rect 16316 11450 16340 11452
rect 16396 11450 16420 11452
rect 16476 11450 16500 11452
rect 16236 11398 16246 11450
rect 16490 11398 16500 11450
rect 16236 11396 16260 11398
rect 16316 11396 16340 11398
rect 16396 11396 16420 11398
rect 16476 11396 16500 11398
rect 16180 11387 16556 11396
rect 16776 11150 16804 11766
rect 17236 11150 17264 11852
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11354 17356 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 11234 17448 12242
rect 17328 11206 17448 11234
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 16028 11076 16080 11082
rect 16028 11018 16080 11024
rect 16920 10908 17296 10917
rect 16976 10906 17000 10908
rect 17056 10906 17080 10908
rect 17136 10906 17160 10908
rect 17216 10906 17240 10908
rect 16976 10854 16986 10906
rect 17230 10854 17240 10906
rect 16976 10852 17000 10854
rect 17056 10852 17080 10854
rect 17136 10852 17160 10854
rect 17216 10852 17240 10854
rect 16920 10843 17296 10852
rect 16180 10364 16556 10373
rect 16236 10362 16260 10364
rect 16316 10362 16340 10364
rect 16396 10362 16420 10364
rect 16476 10362 16500 10364
rect 16236 10310 16246 10362
rect 16490 10310 16500 10362
rect 16236 10308 16260 10310
rect 16316 10308 16340 10310
rect 16396 10308 16420 10310
rect 16476 10308 16500 10310
rect 16180 10299 16556 10308
rect 16920 9820 17296 9829
rect 16976 9818 17000 9820
rect 17056 9818 17080 9820
rect 17136 9818 17160 9820
rect 17216 9818 17240 9820
rect 16976 9766 16986 9818
rect 17230 9766 17240 9818
rect 16976 9764 17000 9766
rect 17056 9764 17080 9766
rect 17136 9764 17160 9766
rect 17216 9764 17240 9766
rect 16920 9755 17296 9764
rect 17328 9518 17356 11206
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17420 9722 17448 9862
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8022 15976 8910
rect 16040 8838 16068 9318
rect 16180 9276 16556 9285
rect 16236 9274 16260 9276
rect 16316 9274 16340 9276
rect 16396 9274 16420 9276
rect 16476 9274 16500 9276
rect 16236 9222 16246 9274
rect 16490 9222 16500 9274
rect 16236 9220 16260 9222
rect 16316 9220 16340 9222
rect 16396 9220 16420 9222
rect 16476 9220 16500 9222
rect 16180 9211 16556 9220
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16592 8498 16620 9318
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16488 8424 16540 8430
rect 16540 8372 16620 8378
rect 16488 8366 16620 8372
rect 16500 8350 16620 8366
rect 16684 8362 16712 8842
rect 16920 8732 17296 8741
rect 16976 8730 17000 8732
rect 17056 8730 17080 8732
rect 17136 8730 17160 8732
rect 17216 8730 17240 8732
rect 16976 8678 16986 8730
rect 17230 8678 17240 8730
rect 16976 8676 17000 8678
rect 17056 8676 17080 8678
rect 17136 8676 17160 8678
rect 17216 8676 17240 8678
rect 16920 8667 17296 8676
rect 16592 8242 16620 8350
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16592 8214 16712 8242
rect 16180 8188 16556 8197
rect 16236 8186 16260 8188
rect 16316 8186 16340 8188
rect 16396 8186 16420 8188
rect 16476 8186 16500 8188
rect 16236 8134 16246 8186
rect 16490 8134 16500 8186
rect 16236 8132 16260 8134
rect 16316 8132 16340 8134
rect 16396 8132 16420 8134
rect 16476 8132 16500 8134
rect 16180 8123 16556 8132
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 16684 7750 16712 8214
rect 17328 7954 17356 9454
rect 17512 8906 17540 12718
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17604 12238 17632 12582
rect 17696 12306 17724 17054
rect 17788 12782 17816 18158
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17202 17908 17478
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17868 15428 17920 15434
rect 17868 15370 17920 15376
rect 17880 14958 17908 15370
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17972 14890 18000 17614
rect 18156 17202 18184 31758
rect 18800 31754 18828 31894
rect 29656 31822 29684 33796
rect 18880 31816 18932 31822
rect 24492 31816 24544 31822
rect 18880 31758 18932 31764
rect 24490 31784 24492 31793
rect 29644 31816 29696 31822
rect 24544 31784 24546 31793
rect 18708 31726 18828 31754
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 18340 31482 18368 31622
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18708 31278 18736 31726
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30394 18736 31214
rect 18696 30388 18748 30394
rect 18696 30330 18748 30336
rect 18708 26382 18736 30330
rect 18892 30122 18920 31758
rect 29644 31758 29696 31764
rect 24490 31719 24546 31728
rect 26700 31680 26752 31686
rect 26700 31622 26752 31628
rect 22920 31580 23296 31589
rect 22976 31578 23000 31580
rect 23056 31578 23080 31580
rect 23136 31578 23160 31580
rect 23216 31578 23240 31580
rect 22976 31526 22986 31578
rect 23230 31526 23240 31578
rect 22976 31524 23000 31526
rect 23056 31524 23080 31526
rect 23136 31524 23160 31526
rect 23216 31524 23240 31526
rect 22920 31515 23296 31524
rect 21088 31408 21140 31414
rect 21088 31350 21140 31356
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 19800 31272 19852 31278
rect 19800 31214 19852 31220
rect 19812 30938 19840 31214
rect 20536 31136 20588 31142
rect 20536 31078 20588 31084
rect 19800 30932 19852 30938
rect 19800 30874 19852 30880
rect 18880 30116 18932 30122
rect 18880 30058 18932 30064
rect 18892 29646 18920 30058
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19616 29572 19668 29578
rect 19616 29514 19668 29520
rect 19352 29102 19380 29514
rect 19628 29238 19656 29514
rect 19812 29306 19840 30874
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19996 30326 20024 30670
rect 20548 30666 20576 31078
rect 20536 30660 20588 30666
rect 20536 30602 20588 30608
rect 20732 30394 20760 31282
rect 21100 30666 21128 31350
rect 21364 31340 21416 31346
rect 21364 31282 21416 31288
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 21088 30660 21140 30666
rect 21088 30602 21140 30608
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19892 29640 19944 29646
rect 19892 29582 19944 29588
rect 19800 29300 19852 29306
rect 19800 29242 19852 29248
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19616 29232 19668 29238
rect 19616 29174 19668 29180
rect 18880 29096 18932 29102
rect 18880 29038 18932 29044
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 18892 28626 18920 29038
rect 18880 28620 18932 28626
rect 18880 28562 18932 28568
rect 18696 26376 18748 26382
rect 18694 26344 18696 26353
rect 18748 26344 18750 26353
rect 18694 26279 18750 26288
rect 18892 25362 18920 28562
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19260 28218 19288 28358
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 19352 27946 19380 29038
rect 19340 27940 19392 27946
rect 19340 27882 19392 27888
rect 19444 27470 19472 29174
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 23866 18368 25094
rect 18432 24954 18460 25162
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18432 24410 18460 24550
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18892 23526 18920 25298
rect 19628 24886 19656 29174
rect 19904 29170 19932 29582
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19812 28762 19840 29106
rect 19996 29102 20024 30262
rect 21100 30258 21128 30602
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 21376 30054 21404 31282
rect 21640 31272 21692 31278
rect 21640 31214 21692 31220
rect 23296 31272 23348 31278
rect 23296 31214 23348 31220
rect 21548 31136 21600 31142
rect 21548 31078 21600 31084
rect 21560 30938 21588 31078
rect 21548 30932 21600 30938
rect 21548 30874 21600 30880
rect 21652 30598 21680 31214
rect 21824 31136 21876 31142
rect 21824 31078 21876 31084
rect 22744 31136 22796 31142
rect 22744 31078 22796 31084
rect 21640 30592 21692 30598
rect 21640 30534 21692 30540
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 21364 30048 21416 30054
rect 21364 29990 21416 29996
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20824 29306 20852 29446
rect 20720 29300 20772 29306
rect 20720 29242 20772 29248
rect 20812 29300 20864 29306
rect 20812 29242 20864 29248
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 19800 28756 19852 28762
rect 19800 28698 19852 28704
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19720 27334 19748 28358
rect 19708 27328 19760 27334
rect 19708 27270 19760 27276
rect 19720 26586 19748 27270
rect 19996 26926 20024 29038
rect 20364 28558 20392 29106
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19996 26382 20024 26862
rect 20260 26512 20312 26518
rect 20260 26454 20312 26460
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19996 25974 20024 26318
rect 19984 25968 20036 25974
rect 19984 25910 20036 25916
rect 20272 25838 20300 26454
rect 20260 25832 20312 25838
rect 20260 25774 20312 25780
rect 19800 25288 19852 25294
rect 19800 25230 19852 25236
rect 19616 24880 19668 24886
rect 19616 24822 19668 24828
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 19338 23488 19394 23497
rect 18328 22432 18380 22438
rect 18328 22374 18380 22380
rect 18340 20874 18368 22374
rect 18892 22098 18920 23462
rect 19338 23423 19394 23432
rect 19352 23118 19380 23423
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18880 22092 18932 22098
rect 19628 22094 19656 24822
rect 19812 24750 19840 25230
rect 20364 24818 20392 28494
rect 20732 27878 20760 29242
rect 20916 28626 20944 29990
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 21008 28762 21036 29582
rect 20996 28756 21048 28762
rect 20996 28698 21048 28704
rect 20904 28620 20956 28626
rect 20904 28562 20956 28568
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 20456 27130 20484 27270
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19904 24410 19932 24618
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 19892 24404 19944 24410
rect 19892 24346 19944 24352
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19996 23730 20024 24074
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 20180 22094 20208 24346
rect 20272 23866 20300 24550
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20260 23520 20312 23526
rect 20260 23462 20312 23468
rect 18880 22034 18932 22040
rect 19444 22066 19656 22094
rect 19444 21962 19472 22066
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19352 21049 19380 21082
rect 19338 21040 19394 21049
rect 19628 21010 19656 22066
rect 19996 22066 20208 22094
rect 19800 21956 19852 21962
rect 19800 21898 19852 21904
rect 19338 20975 19394 20984
rect 19616 21004 19668 21010
rect 19616 20946 19668 20952
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18248 19242 18276 20810
rect 18236 19236 18288 19242
rect 18236 19178 18288 19184
rect 18248 18873 18276 19178
rect 18234 18864 18290 18873
rect 18234 18799 18290 18808
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16794 18092 16934
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18156 16250 18184 17138
rect 18248 16402 18276 17546
rect 18340 17218 18368 20810
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18616 19854 18644 20470
rect 19076 19990 19104 20810
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 18604 19848 18656 19854
rect 18524 19808 18604 19836
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 18432 17338 18460 18294
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18340 17190 18460 17218
rect 18432 17134 18460 17190
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18432 16658 18460 17070
rect 18420 16652 18472 16658
rect 18420 16594 18472 16600
rect 18248 16374 18460 16402
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18340 16130 18368 16186
rect 18248 16114 18368 16130
rect 18236 16108 18368 16114
rect 18288 16102 18368 16108
rect 18236 16050 18288 16056
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18340 15502 18368 15642
rect 18328 15496 18380 15502
rect 18328 15438 18380 15444
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 15162 18092 15302
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17880 14074 17908 14282
rect 17972 14278 18000 14826
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17880 11286 17908 12038
rect 18064 11762 18092 12038
rect 18156 11898 18184 12718
rect 18144 11892 18196 11898
rect 18196 11852 18276 11880
rect 18144 11834 18196 11840
rect 18248 11762 18276 11852
rect 18340 11762 18368 13194
rect 18432 12306 18460 16374
rect 18524 16250 18552 19808
rect 18604 19790 18656 19796
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18604 19236 18656 19242
rect 18604 19178 18656 19184
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 15434 18552 15982
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18524 14958 18552 15370
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18524 14618 18552 14894
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18616 13258 18644 19178
rect 18892 19174 18920 19654
rect 19168 19514 19196 19926
rect 19260 19718 19288 20470
rect 19708 20256 19760 20262
rect 19708 20198 19760 20204
rect 19340 19984 19392 19990
rect 19392 19944 19564 19972
rect 19340 19926 19392 19932
rect 19340 19848 19392 19854
rect 19338 19816 19340 19825
rect 19432 19848 19484 19854
rect 19392 19816 19394 19825
rect 19484 19802 19491 19836
rect 19536 19802 19564 19944
rect 19484 19796 19564 19802
rect 19432 19790 19564 19796
rect 19463 19774 19564 19790
rect 19338 19751 19394 19760
rect 19248 19712 19300 19718
rect 19720 19666 19748 20198
rect 19248 19654 19300 19660
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19260 19446 19288 19654
rect 19463 19638 19748 19666
rect 19463 19530 19491 19638
rect 19812 19530 19840 21898
rect 19996 21146 20024 22066
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20180 21146 20208 21898
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20088 19961 20116 20878
rect 20074 19952 20130 19961
rect 20074 19887 20130 19896
rect 19892 19848 19944 19854
rect 19890 19816 19892 19825
rect 19944 19816 19946 19825
rect 20272 19786 20300 23462
rect 20364 21706 20392 24754
rect 20456 24206 20484 26318
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24206 20668 25094
rect 20824 24818 20852 25162
rect 20812 24812 20864 24818
rect 20812 24754 20864 24760
rect 20916 24750 20944 28562
rect 21652 28082 21680 30534
rect 21836 30394 21864 31078
rect 22180 31036 22556 31045
rect 22236 31034 22260 31036
rect 22316 31034 22340 31036
rect 22396 31034 22420 31036
rect 22476 31034 22500 31036
rect 22236 30982 22246 31034
rect 22490 30982 22500 31034
rect 22236 30980 22260 30982
rect 22316 30980 22340 30982
rect 22396 30980 22420 30982
rect 22476 30980 22500 30982
rect 22180 30971 22556 30980
rect 22756 30394 22784 31078
rect 23308 30938 23336 31214
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 24124 31136 24176 31142
rect 24124 31078 24176 31084
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 21824 30388 21876 30394
rect 21824 30330 21876 30336
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 21916 29776 21968 29782
rect 21916 29718 21968 29724
rect 21824 28960 21876 28966
rect 21824 28902 21876 28908
rect 21836 28558 21864 28902
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21640 28076 21692 28082
rect 21640 28018 21692 28024
rect 21928 27962 21956 29718
rect 22112 28422 22140 30194
rect 22180 29948 22556 29957
rect 22236 29946 22260 29948
rect 22316 29946 22340 29948
rect 22396 29946 22420 29948
rect 22476 29946 22500 29948
rect 22236 29894 22246 29946
rect 22490 29894 22500 29946
rect 22236 29892 22260 29894
rect 22316 29892 22340 29894
rect 22396 29892 22420 29894
rect 22476 29892 22500 29894
rect 22180 29883 22556 29892
rect 22848 29646 22876 30874
rect 24044 30666 24072 31078
rect 24136 30938 24164 31078
rect 24228 30938 24256 31282
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24688 30938 24716 31214
rect 24124 30932 24176 30938
rect 24124 30874 24176 30880
rect 24216 30932 24268 30938
rect 24216 30874 24268 30880
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 23664 30660 23716 30666
rect 23664 30602 23716 30608
rect 24032 30660 24084 30666
rect 24032 30602 24084 30608
rect 22920 30492 23296 30501
rect 22976 30490 23000 30492
rect 23056 30490 23080 30492
rect 23136 30490 23160 30492
rect 23216 30490 23240 30492
rect 22976 30438 22986 30490
rect 23230 30438 23240 30490
rect 22976 30436 23000 30438
rect 23056 30436 23080 30438
rect 23136 30436 23160 30438
rect 23216 30436 23240 30438
rect 22920 30427 23296 30436
rect 23676 30274 23704 30602
rect 23216 30258 23704 30274
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23204 30252 23704 30258
rect 23256 30246 23704 30252
rect 23204 30194 23256 30200
rect 23032 29850 23060 30194
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23020 29844 23072 29850
rect 23020 29786 23072 29792
rect 23124 29646 23152 29990
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23388 29504 23440 29510
rect 23388 29446 23440 29452
rect 22920 29404 23296 29413
rect 22976 29402 23000 29404
rect 23056 29402 23080 29404
rect 23136 29402 23160 29404
rect 23216 29402 23240 29404
rect 22976 29350 22986 29402
rect 23230 29350 23240 29402
rect 22976 29348 23000 29350
rect 23056 29348 23080 29350
rect 23136 29348 23160 29350
rect 23216 29348 23240 29350
rect 22920 29339 23296 29348
rect 22836 29096 22888 29102
rect 22836 29038 22888 29044
rect 22180 28860 22556 28869
rect 22236 28858 22260 28860
rect 22316 28858 22340 28860
rect 22396 28858 22420 28860
rect 22476 28858 22500 28860
rect 22236 28806 22246 28858
rect 22490 28806 22500 28858
rect 22236 28804 22260 28806
rect 22316 28804 22340 28806
rect 22396 28804 22420 28806
rect 22476 28804 22500 28806
rect 22180 28795 22556 28804
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 22284 28144 22336 28150
rect 22204 28092 22284 28098
rect 22204 28086 22336 28092
rect 22204 28070 22324 28086
rect 22468 28076 22520 28082
rect 22204 27962 22232 28070
rect 22468 28018 22520 28024
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22480 27985 22508 28018
rect 21824 27940 21876 27946
rect 21928 27934 22232 27962
rect 22466 27976 22522 27985
rect 22466 27911 22522 27920
rect 21824 27882 21876 27888
rect 20996 27532 21048 27538
rect 20996 27474 21048 27480
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20456 23186 20484 24142
rect 20444 23180 20496 23186
rect 20496 23140 20576 23168
rect 20444 23122 20496 23128
rect 20548 22098 20576 23140
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 20364 21690 20760 21706
rect 20352 21684 20760 21690
rect 20404 21678 20760 21684
rect 20352 21626 20404 21632
rect 20732 20534 20760 21678
rect 20916 21486 20944 24686
rect 21008 24274 21036 27474
rect 21548 27464 21600 27470
rect 21836 27452 21864 27882
rect 22180 27772 22556 27781
rect 22236 27770 22260 27772
rect 22316 27770 22340 27772
rect 22396 27770 22420 27772
rect 22476 27770 22500 27772
rect 22236 27718 22246 27770
rect 22490 27718 22500 27770
rect 22236 27716 22260 27718
rect 22316 27716 22340 27718
rect 22396 27716 22420 27718
rect 22476 27716 22500 27718
rect 22180 27707 22556 27716
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 21916 27464 21968 27470
rect 21836 27424 21916 27452
rect 21548 27406 21600 27412
rect 21916 27406 21968 27412
rect 21560 27130 21588 27406
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21376 26314 21404 26726
rect 21836 26586 21864 26862
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 21364 26308 21416 26314
rect 21364 26250 21416 26256
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 20996 24268 21048 24274
rect 20996 24210 21048 24216
rect 21008 23526 21036 24210
rect 21192 23866 21220 24550
rect 21284 24410 21312 24686
rect 21376 24410 21404 24754
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21284 23118 21312 24346
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23866 21864 24006
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21928 23746 21956 27406
rect 22020 27130 22048 27610
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 22388 27130 22416 27542
rect 22664 27538 22692 28018
rect 22848 27554 22876 29038
rect 22920 28316 23296 28325
rect 22976 28314 23000 28316
rect 23056 28314 23080 28316
rect 23136 28314 23160 28316
rect 23216 28314 23240 28316
rect 22976 28262 22986 28314
rect 23230 28262 23240 28314
rect 22976 28260 23000 28262
rect 23056 28260 23080 28262
rect 23136 28260 23160 28262
rect 23216 28260 23240 28262
rect 22920 28251 23296 28260
rect 23400 28082 23428 29446
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 22940 27674 22968 28018
rect 23386 27976 23442 27985
rect 23386 27911 23442 27920
rect 23480 27940 23532 27946
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 22848 27538 22968 27554
rect 22652 27532 22704 27538
rect 22848 27532 22980 27538
rect 22848 27526 22928 27532
rect 22652 27474 22704 27480
rect 22928 27474 22980 27480
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 22376 27124 22428 27130
rect 22376 27066 22428 27072
rect 22480 27062 22508 27270
rect 22468 27056 22520 27062
rect 22468 26998 22520 27004
rect 22572 26926 22600 27270
rect 22560 26920 22612 26926
rect 22560 26862 22612 26868
rect 22664 26858 22692 27474
rect 23032 27384 23060 27814
rect 23400 27470 23428 27911
rect 23480 27882 23532 27888
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 22756 27356 23060 27384
rect 22652 26852 22704 26858
rect 22652 26794 22704 26800
rect 22180 26684 22556 26693
rect 22236 26682 22260 26684
rect 22316 26682 22340 26684
rect 22396 26682 22420 26684
rect 22476 26682 22500 26684
rect 22236 26630 22246 26682
rect 22490 26630 22500 26682
rect 22236 26628 22260 26630
rect 22316 26628 22340 26630
rect 22396 26628 22420 26630
rect 22476 26628 22500 26630
rect 22180 26619 22556 26628
rect 22180 25596 22556 25605
rect 22236 25594 22260 25596
rect 22316 25594 22340 25596
rect 22396 25594 22420 25596
rect 22476 25594 22500 25596
rect 22236 25542 22246 25594
rect 22490 25542 22500 25594
rect 22236 25540 22260 25542
rect 22316 25540 22340 25542
rect 22396 25540 22420 25542
rect 22476 25540 22500 25542
rect 22180 25531 22556 25540
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22112 24342 22140 24550
rect 22180 24508 22556 24517
rect 22236 24506 22260 24508
rect 22316 24506 22340 24508
rect 22396 24506 22420 24508
rect 22476 24506 22500 24508
rect 22236 24454 22246 24506
rect 22490 24454 22500 24506
rect 22236 24452 22260 24454
rect 22316 24452 22340 24454
rect 22396 24452 22420 24454
rect 22476 24452 22500 24454
rect 22180 24443 22556 24452
rect 22100 24336 22152 24342
rect 22100 24278 22152 24284
rect 21836 23718 21956 23746
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21836 22982 21864 23718
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22112 23118 22140 23530
rect 22180 23420 22556 23429
rect 22236 23418 22260 23420
rect 22316 23418 22340 23420
rect 22396 23418 22420 23420
rect 22476 23418 22500 23420
rect 22236 23366 22246 23418
rect 22490 23366 22500 23418
rect 22236 23364 22260 23366
rect 22316 23364 22340 23366
rect 22396 23364 22420 23366
rect 22476 23364 22500 23366
rect 22180 23355 22556 23364
rect 22664 23322 22692 23734
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 20994 21992 21050 22001
rect 20994 21927 21050 21936
rect 21008 21894 21036 21927
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21836 21622 21864 22918
rect 22180 22332 22556 22341
rect 22236 22330 22260 22332
rect 22316 22330 22340 22332
rect 22396 22330 22420 22332
rect 22476 22330 22500 22332
rect 22236 22278 22246 22330
rect 22490 22278 22500 22330
rect 22236 22276 22260 22278
rect 22316 22276 22340 22278
rect 22396 22276 22420 22278
rect 22476 22276 22500 22278
rect 22180 22267 22556 22276
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 22112 21146 22140 21490
rect 22180 21244 22556 21253
rect 22236 21242 22260 21244
rect 22316 21242 22340 21244
rect 22396 21242 22420 21244
rect 22476 21242 22500 21244
rect 22236 21190 22246 21242
rect 22490 21190 22500 21242
rect 22236 21188 22260 21190
rect 22316 21188 22340 21190
rect 22396 21188 22420 21190
rect 22476 21188 22500 21190
rect 22180 21179 22556 21188
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 21652 20998 21956 21026
rect 21652 20942 21680 20998
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21008 20534 21036 20878
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20812 20324 20864 20330
rect 20812 20266 20864 20272
rect 20824 19854 20852 20266
rect 20916 19922 20944 20334
rect 21376 19938 21404 20402
rect 21376 19922 21496 19938
rect 20904 19916 20956 19922
rect 21376 19916 21508 19922
rect 21376 19910 21456 19916
rect 20904 19858 20956 19864
rect 21456 19858 21508 19864
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 19890 19751 19946 19760
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 19444 19502 19491 19530
rect 19536 19502 19840 19530
rect 19248 19440 19300 19446
rect 19248 19382 19300 19388
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 19260 18290 19288 19382
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 18694 17776 18750 17785
rect 18694 17711 18696 17720
rect 18748 17711 18750 17720
rect 18696 17682 18748 17688
rect 18984 17542 19012 18226
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17134 19012 17478
rect 19076 17270 19104 17614
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18708 15978 18736 16526
rect 18788 16448 18840 16454
rect 18984 16436 19012 17070
rect 19076 16794 19104 17070
rect 19064 16788 19116 16794
rect 19064 16730 19116 16736
rect 19168 16538 19196 17614
rect 19260 17202 19288 17818
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 19352 17649 19380 17682
rect 19444 17678 19472 19502
rect 19432 17672 19484 17678
rect 19338 17640 19394 17649
rect 19432 17614 19484 17620
rect 19338 17575 19394 17584
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19260 16658 19288 17138
rect 19444 16794 19472 17614
rect 19536 17338 19564 19502
rect 20456 19378 20484 19722
rect 20626 19408 20682 19417
rect 19616 19372 19668 19378
rect 20444 19372 20496 19378
rect 19668 19320 19932 19334
rect 19616 19314 19932 19320
rect 20626 19343 20682 19352
rect 20444 19314 20496 19320
rect 19628 19306 19932 19314
rect 20640 19310 20668 19343
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19720 18290 19748 18702
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19628 17542 19656 18090
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19168 16522 19288 16538
rect 19168 16516 19300 16522
rect 19168 16510 19248 16516
rect 19248 16458 19300 16464
rect 19156 16448 19208 16454
rect 18984 16408 19156 16436
rect 18788 16390 18840 16396
rect 19156 16390 19208 16396
rect 18800 16250 18828 16390
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 19168 16114 19196 16390
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18708 14006 18736 15914
rect 19168 15706 19196 16050
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19260 15434 19288 16458
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19352 14822 19380 16390
rect 19444 15706 19472 16730
rect 19614 16280 19670 16289
rect 19614 16215 19670 16224
rect 19628 16114 19656 16215
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19628 15978 19656 16050
rect 19616 15972 19668 15978
rect 19616 15914 19668 15920
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19720 15502 19748 18226
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18616 11762 18644 12922
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12238 18736 12582
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18340 11354 18368 11698
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17866 8800 17922 8809
rect 17866 8735 17922 8744
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17880 7750 17908 8735
rect 17972 8498 18000 8910
rect 18064 8838 18092 9998
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18248 8906 18276 9386
rect 18340 8974 18368 9590
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18236 8900 18288 8906
rect 18236 8842 18288 8848
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18616 8498 18644 11698
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18708 8566 18736 11290
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8566 18828 8774
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 16316 7546 16344 7686
rect 16920 7644 17296 7653
rect 16976 7642 17000 7644
rect 17056 7642 17080 7644
rect 17136 7642 17160 7644
rect 17216 7642 17240 7644
rect 16976 7590 16986 7642
rect 17230 7590 17240 7642
rect 16976 7588 17000 7590
rect 17056 7588 17080 7590
rect 17136 7588 17160 7590
rect 17216 7588 17240 7590
rect 16920 7579 17296 7588
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16180 7100 16556 7109
rect 16236 7098 16260 7100
rect 16316 7098 16340 7100
rect 16396 7098 16420 7100
rect 16476 7098 16500 7100
rect 16236 7046 16246 7098
rect 16490 7046 16500 7098
rect 16236 7044 16260 7046
rect 16316 7044 16340 7046
rect 16396 7044 16420 7046
rect 16476 7044 16500 7046
rect 16180 7035 16556 7044
rect 16920 6556 17296 6565
rect 16976 6554 17000 6556
rect 17056 6554 17080 6556
rect 17136 6554 17160 6556
rect 17216 6554 17240 6556
rect 16976 6502 16986 6554
rect 17230 6502 17240 6554
rect 16976 6500 17000 6502
rect 17056 6500 17080 6502
rect 17136 6500 17160 6502
rect 17216 6500 17240 6502
rect 16920 6491 17296 6500
rect 17972 6322 18000 8434
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18340 6798 18368 7958
rect 18616 7886 18644 8434
rect 18708 7886 18736 8502
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 16180 6012 16556 6021
rect 16236 6010 16260 6012
rect 16316 6010 16340 6012
rect 16396 6010 16420 6012
rect 16476 6010 16500 6012
rect 16236 5958 16246 6010
rect 16490 5958 16500 6010
rect 16236 5956 16260 5958
rect 16316 5956 16340 5958
rect 16396 5956 16420 5958
rect 16476 5956 16500 5958
rect 16180 5947 16556 5956
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 16920 5468 17296 5477
rect 16976 5466 17000 5468
rect 17056 5466 17080 5468
rect 17136 5466 17160 5468
rect 17216 5466 17240 5468
rect 16976 5414 16986 5466
rect 17230 5414 17240 5466
rect 16976 5412 17000 5414
rect 17056 5412 17080 5414
rect 17136 5412 17160 5414
rect 17216 5412 17240 5414
rect 16920 5403 17296 5412
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 16180 4924 16556 4933
rect 16236 4922 16260 4924
rect 16316 4922 16340 4924
rect 16396 4922 16420 4924
rect 16476 4922 16500 4924
rect 16236 4870 16246 4922
rect 16490 4870 16500 4922
rect 16236 4868 16260 4870
rect 16316 4868 16340 4870
rect 16396 4868 16420 4870
rect 16476 4868 16500 4870
rect 16180 4859 16556 4868
rect 15856 4814 16068 4842
rect 15936 4752 15988 4758
rect 15764 4700 15936 4706
rect 15764 4694 15988 4700
rect 15764 4678 15976 4694
rect 16040 4690 16068 4814
rect 16592 4690 16620 4966
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 17420 4622 17448 4966
rect 17788 4622 17816 5238
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 14936 4214 14964 4422
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14844 3602 14872 4014
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13924 2446 13952 3538
rect 15396 3398 15424 3878
rect 15948 3466 15976 4422
rect 16684 4282 16712 4422
rect 16920 4380 17296 4389
rect 16976 4378 17000 4380
rect 17056 4378 17080 4380
rect 17136 4378 17160 4380
rect 17216 4378 17240 4380
rect 16976 4326 16986 4378
rect 17230 4326 17240 4378
rect 16976 4324 17000 4326
rect 17056 4324 17080 4326
rect 17136 4324 17160 4326
rect 17216 4324 17240 4326
rect 16920 4315 17296 4324
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 17696 4146 17724 4558
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 4146 18000 4422
rect 18432 4282 18460 4490
rect 18420 4276 18472 4282
rect 18420 4218 18472 4224
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 16180 3836 16556 3845
rect 16236 3834 16260 3836
rect 16316 3834 16340 3836
rect 16396 3834 16420 3836
rect 16476 3834 16500 3836
rect 16236 3782 16246 3834
rect 16490 3782 16500 3834
rect 16236 3780 16260 3782
rect 16316 3780 16340 3782
rect 16396 3780 16420 3782
rect 16476 3780 16500 3782
rect 16180 3771 16556 3780
rect 17144 3738 17172 4082
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17696 3602 17724 3878
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 16920 3292 17296 3301
rect 16976 3290 17000 3292
rect 17056 3290 17080 3292
rect 17136 3290 17160 3292
rect 17216 3290 17240 3292
rect 16976 3238 16986 3290
rect 17230 3238 17240 3290
rect 16976 3236 17000 3238
rect 17056 3236 17080 3238
rect 17136 3236 17160 3238
rect 17216 3236 17240 3238
rect 16920 3227 17296 3236
rect 18984 2774 19012 14758
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19444 12986 19472 13194
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19076 11898 19104 12786
rect 19340 12164 19392 12170
rect 19340 12106 19392 12112
rect 19352 11914 19380 12106
rect 19444 12102 19472 12922
rect 19720 12714 19748 15438
rect 19812 12782 19840 18906
rect 19904 17882 19932 19306
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20732 18222 20760 19722
rect 20916 19378 20944 19858
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21008 19378 21036 19790
rect 21560 19786 21588 20538
rect 21652 20380 21680 20742
rect 21744 20602 21772 20878
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21732 20392 21784 20398
rect 21652 20352 21732 20380
rect 21732 20334 21784 20340
rect 21744 19854 21772 20334
rect 21836 19990 21864 20538
rect 21928 20466 21956 20998
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20602 22232 20742
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22112 20058 22140 20334
rect 22480 20262 22508 20946
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22572 20466 22600 20742
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22180 20156 22556 20165
rect 22236 20154 22260 20156
rect 22316 20154 22340 20156
rect 22396 20154 22420 20156
rect 22476 20154 22500 20156
rect 22236 20102 22246 20154
rect 22490 20102 22500 20154
rect 22236 20100 22260 20102
rect 22316 20100 22340 20102
rect 22396 20100 22420 20102
rect 22476 20100 22500 20102
rect 22180 20091 22556 20100
rect 22664 20058 22692 23054
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22652 20052 22704 20058
rect 22652 19994 22704 20000
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21548 19780 21600 19786
rect 21548 19722 21600 19728
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 19378 21128 19654
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20076 18080 20128 18086
rect 20076 18022 20128 18028
rect 19892 17876 19944 17882
rect 19892 17818 19944 17824
rect 20088 17678 20116 18022
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19904 16454 19932 17614
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20272 17338 20300 17546
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20916 17134 20944 19314
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 21008 17066 21036 19314
rect 21284 19310 21312 19722
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 19446 21496 19654
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21086 17640 21142 17649
rect 21086 17575 21142 17584
rect 21100 17542 21128 17575
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16794 20760 16934
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 19892 16448 19944 16454
rect 19892 16390 19944 16396
rect 20088 16114 20116 16458
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16289 21036 16390
rect 20994 16280 21050 16289
rect 20994 16215 21050 16224
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20916 15570 20944 16050
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 15026 20576 15302
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 13462 20668 14758
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 21100 12986 21128 17478
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19708 12708 19760 12714
rect 19708 12650 19760 12656
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19064 11892 19116 11898
rect 19352 11886 19472 11914
rect 19064 11834 19116 11840
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19352 10826 19380 11018
rect 19260 10798 19380 10826
rect 19260 9654 19288 10798
rect 19444 10130 19472 11886
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19064 9512 19116 9518
rect 19064 9454 19116 9460
rect 19076 8634 19104 9454
rect 19168 9178 19196 9522
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19260 9178 19288 9454
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 19156 8968 19208 8974
rect 19352 8956 19380 9862
rect 19628 9178 19656 9862
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19208 8928 19380 8956
rect 19156 8910 19208 8916
rect 19628 8634 19656 9114
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19812 8430 19840 12718
rect 20364 12434 20392 12786
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20640 12442 20668 12718
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12436 20680 12442
rect 20364 12406 20484 12434
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 11218 20392 11698
rect 20456 11626 20484 12406
rect 20628 12378 20680 12384
rect 20732 12220 20760 12582
rect 20904 12232 20956 12238
rect 20732 12192 20904 12220
rect 20904 12174 20956 12180
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11762 21036 12038
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 8634 19932 9522
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19812 6866 19840 8366
rect 19800 6860 19852 6866
rect 19800 6802 19852 6808
rect 19432 6792 19484 6798
rect 19484 6740 19840 6746
rect 19432 6734 19840 6740
rect 19444 6718 19840 6734
rect 19812 6662 19840 6718
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19168 6338 19196 6598
rect 19260 6458 19288 6598
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19168 6310 19380 6338
rect 19352 6118 19380 6310
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19720 5574 19748 6598
rect 19996 5778 20024 10066
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20824 9586 20852 9998
rect 21100 9674 21128 12922
rect 21192 12850 21220 19246
rect 21284 18698 21312 19246
rect 21560 19174 21588 19722
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21560 18766 21588 19110
rect 21652 18834 21680 19722
rect 21744 18970 21772 19790
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21916 19712 21968 19718
rect 21916 19654 21968 19660
rect 21732 18964 21784 18970
rect 21732 18906 21784 18912
rect 21836 18902 21864 19654
rect 21928 19310 21956 19654
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 21272 18692 21324 18698
rect 21272 18634 21324 18640
rect 21284 18086 21312 18634
rect 21560 18290 21588 18702
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21284 17134 21312 18022
rect 21376 17678 21404 18022
rect 21836 17678 21864 18566
rect 22112 17678 22140 19314
rect 22572 19156 22600 19450
rect 22664 19378 22692 19790
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22572 19128 22692 19156
rect 22180 19068 22556 19077
rect 22236 19066 22260 19068
rect 22316 19066 22340 19068
rect 22396 19066 22420 19068
rect 22476 19066 22500 19068
rect 22236 19014 22246 19066
rect 22490 19014 22500 19066
rect 22236 19012 22260 19014
rect 22316 19012 22340 19014
rect 22396 19012 22420 19014
rect 22476 19012 22500 19014
rect 22180 19003 22556 19012
rect 22180 17980 22556 17989
rect 22236 17978 22260 17980
rect 22316 17978 22340 17980
rect 22396 17978 22420 17980
rect 22476 17978 22500 17980
rect 22236 17926 22246 17978
rect 22490 17926 22500 17978
rect 22236 17924 22260 17926
rect 22316 17924 22340 17926
rect 22396 17924 22420 17926
rect 22476 17924 22500 17926
rect 22180 17915 22556 17924
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 21376 17270 21404 17614
rect 21732 17604 21784 17610
rect 21732 17546 21784 17552
rect 21364 17264 21416 17270
rect 21364 17206 21416 17212
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21744 16794 21772 17546
rect 22112 17202 22140 17614
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21732 16788 21784 16794
rect 21732 16730 21784 16736
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21376 16250 21404 16458
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 12986 21312 15438
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 12986 21404 13670
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21468 12850 21496 13126
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21008 9646 21128 9674
rect 21008 9586 21036 9646
rect 21192 9586 21220 12786
rect 21744 12442 21772 16730
rect 22020 16114 22048 16934
rect 22112 16590 22140 17138
rect 22296 17066 22324 17546
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 17202 22600 17478
rect 22664 17270 22692 19128
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22652 16992 22704 16998
rect 22652 16934 22704 16940
rect 22180 16892 22556 16901
rect 22236 16890 22260 16892
rect 22316 16890 22340 16892
rect 22396 16890 22420 16892
rect 22476 16890 22500 16892
rect 22236 16838 22246 16890
rect 22490 16838 22500 16890
rect 22236 16836 22260 16838
rect 22316 16836 22340 16838
rect 22396 16836 22420 16838
rect 22476 16836 22500 16838
rect 22180 16827 22556 16836
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22112 16182 22140 16526
rect 22100 16176 22152 16182
rect 22100 16118 22152 16124
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22388 16046 22416 16730
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22180 15804 22556 15813
rect 22236 15802 22260 15804
rect 22316 15802 22340 15804
rect 22396 15802 22420 15804
rect 22476 15802 22500 15804
rect 22236 15750 22246 15802
rect 22490 15750 22500 15802
rect 22236 15748 22260 15750
rect 22316 15748 22340 15750
rect 22396 15748 22420 15750
rect 22476 15748 22500 15750
rect 22180 15739 22556 15748
rect 22664 15706 22692 16934
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22020 15162 22048 15370
rect 22008 15156 22060 15162
rect 21928 15116 22008 15144
rect 21928 15026 21956 15116
rect 22008 15098 22060 15104
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14890 22048 14962
rect 22008 14884 22060 14890
rect 22008 14826 22060 14832
rect 22180 14716 22556 14725
rect 22236 14714 22260 14716
rect 22316 14714 22340 14716
rect 22396 14714 22420 14716
rect 22476 14714 22500 14716
rect 22236 14662 22246 14714
rect 22490 14662 22500 14714
rect 22236 14660 22260 14662
rect 22316 14660 22340 14662
rect 22396 14660 22420 14662
rect 22476 14660 22500 14662
rect 22180 14651 22556 14660
rect 22756 14498 22784 27356
rect 22920 27228 23296 27237
rect 22976 27226 23000 27228
rect 23056 27226 23080 27228
rect 23136 27226 23160 27228
rect 23216 27226 23240 27228
rect 22976 27174 22986 27226
rect 23230 27174 23240 27226
rect 22976 27172 23000 27174
rect 23056 27172 23080 27174
rect 23136 27172 23160 27174
rect 23216 27172 23240 27174
rect 22920 27163 23296 27172
rect 23400 27010 23428 27406
rect 23492 27130 23520 27882
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23400 26982 23520 27010
rect 22920 26140 23296 26149
rect 22976 26138 23000 26140
rect 23056 26138 23080 26140
rect 23136 26138 23160 26140
rect 23216 26138 23240 26140
rect 22976 26086 22986 26138
rect 23230 26086 23240 26138
rect 22976 26084 23000 26086
rect 23056 26084 23080 26086
rect 23136 26084 23160 26086
rect 23216 26084 23240 26086
rect 22920 26075 23296 26084
rect 22920 25052 23296 25061
rect 22976 25050 23000 25052
rect 23056 25050 23080 25052
rect 23136 25050 23160 25052
rect 23216 25050 23240 25052
rect 22976 24998 22986 25050
rect 23230 24998 23240 25050
rect 22976 24996 23000 24998
rect 23056 24996 23080 24998
rect 23136 24996 23160 24998
rect 23216 24996 23240 24998
rect 22920 24987 23296 24996
rect 22836 24064 22888 24070
rect 22836 24006 22888 24012
rect 22848 23322 22876 24006
rect 22920 23964 23296 23973
rect 22976 23962 23000 23964
rect 23056 23962 23080 23964
rect 23136 23962 23160 23964
rect 23216 23962 23240 23964
rect 22976 23910 22986 23962
rect 23230 23910 23240 23962
rect 22976 23908 23000 23910
rect 23056 23908 23080 23910
rect 23136 23908 23160 23910
rect 23216 23908 23240 23910
rect 22920 23899 23296 23908
rect 23492 23848 23520 26982
rect 23572 24676 23624 24682
rect 23572 24618 23624 24624
rect 23308 23820 23520 23848
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22836 23316 22888 23322
rect 22836 23258 22888 23264
rect 23032 22964 23060 23462
rect 23124 23118 23152 23462
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23308 23050 23336 23820
rect 23584 23730 23612 24618
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23492 23322 23520 23666
rect 23676 23662 23704 30246
rect 23940 29776 23992 29782
rect 23940 29718 23992 29724
rect 24400 29776 24452 29782
rect 24400 29718 24452 29724
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23768 27130 23796 27950
rect 23756 27124 23808 27130
rect 23756 27066 23808 27072
rect 23860 26790 23888 29446
rect 23848 26784 23900 26790
rect 23848 26726 23900 26732
rect 23848 24608 23900 24614
rect 23848 24550 23900 24556
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 23798 23796 24142
rect 23860 23866 23888 24550
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23756 23792 23808 23798
rect 23756 23734 23808 23740
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23848 23656 23900 23662
rect 23848 23598 23900 23604
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22848 22936 23060 22964
rect 22848 15026 22876 22936
rect 22920 22876 23296 22885
rect 22976 22874 23000 22876
rect 23056 22874 23080 22876
rect 23136 22874 23160 22876
rect 23216 22874 23240 22876
rect 22976 22822 22986 22874
rect 23230 22822 23240 22874
rect 22976 22820 23000 22822
rect 23056 22820 23080 22822
rect 23136 22820 23160 22822
rect 23216 22820 23240 22822
rect 22920 22811 23296 22820
rect 23676 22506 23704 23598
rect 23756 23520 23808 23526
rect 23756 23462 23808 23468
rect 23768 22778 23796 23462
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 22920 21788 23296 21797
rect 22976 21786 23000 21788
rect 23056 21786 23080 21788
rect 23136 21786 23160 21788
rect 23216 21786 23240 21788
rect 22976 21734 22986 21786
rect 23230 21734 23240 21786
rect 22976 21732 23000 21734
rect 23056 21732 23080 21734
rect 23136 21732 23160 21734
rect 23216 21732 23240 21734
rect 22920 21723 23296 21732
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23400 21010 23428 21490
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23492 21010 23520 21422
rect 23768 21146 23796 21966
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 22920 20700 23296 20709
rect 22976 20698 23000 20700
rect 23056 20698 23080 20700
rect 23136 20698 23160 20700
rect 23216 20698 23240 20700
rect 22976 20646 22986 20698
rect 23230 20646 23240 20698
rect 22976 20644 23000 20646
rect 23056 20644 23080 20646
rect 23136 20644 23160 20646
rect 23216 20644 23240 20646
rect 22920 20635 23296 20644
rect 23296 20596 23348 20602
rect 23296 20538 23348 20544
rect 23308 20398 23336 20538
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22940 19990 22968 20198
rect 22928 19984 22980 19990
rect 22928 19926 22980 19932
rect 23124 19854 23152 20334
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23400 19786 23428 20810
rect 23492 20754 23520 20946
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23664 20800 23716 20806
rect 23492 20726 23612 20754
rect 23664 20742 23716 20748
rect 23480 20460 23532 20466
rect 23480 20402 23532 20408
rect 23388 19780 23440 19786
rect 23388 19722 23440 19728
rect 22920 19612 23296 19621
rect 22976 19610 23000 19612
rect 23056 19610 23080 19612
rect 23136 19610 23160 19612
rect 23216 19610 23240 19612
rect 22976 19558 22986 19610
rect 23230 19558 23240 19610
rect 22976 19556 23000 19558
rect 23056 19556 23080 19558
rect 23136 19556 23160 19558
rect 23216 19556 23240 19558
rect 22920 19547 23296 19556
rect 22920 18524 23296 18533
rect 22976 18522 23000 18524
rect 23056 18522 23080 18524
rect 23136 18522 23160 18524
rect 23216 18522 23240 18524
rect 22976 18470 22986 18522
rect 23230 18470 23240 18522
rect 22976 18468 23000 18470
rect 23056 18468 23080 18470
rect 23136 18468 23160 18470
rect 23216 18468 23240 18470
rect 22920 18459 23296 18468
rect 23400 18358 23428 19722
rect 23492 19718 23520 20402
rect 23584 20330 23612 20726
rect 23572 20324 23624 20330
rect 23572 20266 23624 20272
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23584 19530 23612 20266
rect 23676 19854 23704 20742
rect 23768 20534 23796 20878
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23492 19502 23612 19530
rect 23492 19174 23520 19502
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23492 18358 23520 19110
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23584 18358 23612 18838
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 23124 17610 23152 18022
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 22920 17436 23296 17445
rect 22976 17434 23000 17436
rect 23056 17434 23080 17436
rect 23136 17434 23160 17436
rect 23216 17434 23240 17436
rect 22976 17382 22986 17434
rect 23230 17382 23240 17434
rect 22976 17380 23000 17382
rect 23056 17380 23080 17382
rect 23136 17380 23160 17382
rect 23216 17380 23240 17382
rect 22920 17371 23296 17380
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 22940 16590 22968 17138
rect 23400 17134 23428 17682
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23032 16794 23060 17070
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23124 16590 23152 16730
rect 23204 16720 23256 16726
rect 23204 16662 23256 16668
rect 23216 16590 23244 16662
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23204 16584 23256 16590
rect 23256 16532 23428 16538
rect 23204 16526 23428 16532
rect 23216 16510 23428 16526
rect 22920 16348 23296 16357
rect 22976 16346 23000 16348
rect 23056 16346 23080 16348
rect 23136 16346 23160 16348
rect 23216 16346 23240 16348
rect 22976 16294 22986 16346
rect 23230 16294 23240 16346
rect 22976 16292 23000 16294
rect 23056 16292 23080 16294
rect 23136 16292 23160 16294
rect 23216 16292 23240 16294
rect 22920 16283 23296 16292
rect 23400 15978 23428 16510
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 22920 15260 23296 15269
rect 22976 15258 23000 15260
rect 23056 15258 23080 15260
rect 23136 15258 23160 15260
rect 23216 15258 23240 15260
rect 22976 15206 22986 15258
rect 23230 15206 23240 15258
rect 22976 15204 23000 15206
rect 23056 15204 23080 15206
rect 23136 15204 23160 15206
rect 23216 15204 23240 15206
rect 22920 15195 23296 15204
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22756 14470 22876 14498
rect 22180 13628 22556 13637
rect 22236 13626 22260 13628
rect 22316 13626 22340 13628
rect 22396 13626 22420 13628
rect 22476 13626 22500 13628
rect 22236 13574 22246 13626
rect 22490 13574 22500 13626
rect 22236 13572 22260 13574
rect 22316 13572 22340 13574
rect 22396 13572 22420 13574
rect 22476 13572 22500 13574
rect 22180 13563 22556 13572
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21836 12730 21864 12786
rect 21836 12702 21956 12730
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21468 11898 21496 12174
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21744 11898 21772 12106
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21928 11830 21956 12702
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21468 11354 21496 11698
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 21560 11082 21588 11698
rect 21548 11076 21600 11082
rect 21548 11018 21600 11024
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 9722 21956 10406
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20904 9512 20956 9518
rect 20824 9460 20904 9466
rect 20824 9454 20956 9460
rect 20824 9438 20944 9454
rect 20168 8900 20220 8906
rect 20168 8842 20220 8848
rect 20180 8634 20208 8842
rect 20168 8628 20220 8634
rect 20168 8570 20220 8576
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20732 6458 20760 6734
rect 20824 6662 20852 9438
rect 21008 7002 21036 9522
rect 21100 9178 21128 9522
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21100 8634 21128 9114
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21836 8634 21864 8842
rect 22020 8634 22048 9318
rect 22112 8922 22140 13262
rect 22376 13252 22428 13258
rect 22744 13252 22796 13258
rect 22428 13212 22744 13240
rect 22376 13194 22428 13200
rect 22744 13194 22796 13200
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22180 12540 22556 12549
rect 22236 12538 22260 12540
rect 22316 12538 22340 12540
rect 22396 12538 22420 12540
rect 22476 12538 22500 12540
rect 22236 12486 22246 12538
rect 22490 12486 22500 12538
rect 22236 12484 22260 12486
rect 22316 12484 22340 12486
rect 22396 12484 22420 12486
rect 22476 12484 22500 12486
rect 22180 12475 22556 12484
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22180 11452 22556 11461
rect 22236 11450 22260 11452
rect 22316 11450 22340 11452
rect 22396 11450 22420 11452
rect 22476 11450 22500 11452
rect 22236 11398 22246 11450
rect 22490 11398 22500 11450
rect 22236 11396 22260 11398
rect 22316 11396 22340 11398
rect 22396 11396 22420 11398
rect 22476 11396 22500 11398
rect 22180 11387 22556 11396
rect 22664 11286 22692 11494
rect 22652 11280 22704 11286
rect 22652 11222 22704 11228
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 11014 22416 11086
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 22388 10690 22416 10950
rect 22388 10662 22692 10690
rect 22180 10364 22556 10373
rect 22236 10362 22260 10364
rect 22316 10362 22340 10364
rect 22396 10362 22420 10364
rect 22476 10362 22500 10364
rect 22236 10310 22246 10362
rect 22490 10310 22500 10362
rect 22236 10308 22260 10310
rect 22316 10308 22340 10310
rect 22396 10308 22420 10310
rect 22476 10308 22500 10310
rect 22180 10299 22556 10308
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22388 9722 22416 9998
rect 22572 9761 22600 10066
rect 22558 9752 22614 9761
rect 22376 9716 22428 9722
rect 22558 9687 22614 9696
rect 22376 9658 22428 9664
rect 22664 9518 22692 10662
rect 22756 9994 22784 12582
rect 22848 10792 22876 14470
rect 22920 14172 23296 14181
rect 22976 14170 23000 14172
rect 23056 14170 23080 14172
rect 23136 14170 23160 14172
rect 23216 14170 23240 14172
rect 22976 14118 22986 14170
rect 23230 14118 23240 14170
rect 22976 14116 23000 14118
rect 23056 14116 23080 14118
rect 23136 14116 23160 14118
rect 23216 14116 23240 14118
rect 22920 14107 23296 14116
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 22920 13084 23296 13093
rect 22976 13082 23000 13084
rect 23056 13082 23080 13084
rect 23136 13082 23160 13084
rect 23216 13082 23240 13084
rect 22976 13030 22986 13082
rect 23230 13030 23240 13082
rect 22976 13028 23000 13030
rect 23056 13028 23080 13030
rect 23136 13028 23160 13030
rect 23216 13028 23240 13030
rect 22920 13019 23296 13028
rect 23400 12986 23428 13262
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23124 12170 23152 12582
rect 23216 12374 23244 12786
rect 23204 12368 23256 12374
rect 23204 12310 23256 12316
rect 23216 12209 23244 12310
rect 23400 12238 23428 12922
rect 23492 12918 23520 17206
rect 23584 17066 23612 17546
rect 23676 17202 23704 19790
rect 23768 19514 23796 20198
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23860 17354 23888 23598
rect 23952 23066 23980 29718
rect 24308 29504 24360 29510
rect 24308 29446 24360 29452
rect 24320 29034 24348 29446
rect 24412 29170 24440 29718
rect 24492 29708 24544 29714
rect 24492 29650 24544 29656
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 24504 29102 24532 29650
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 29306 24624 29446
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24688 29170 24716 30874
rect 24952 30728 25004 30734
rect 24952 30670 25004 30676
rect 24964 30326 24992 30670
rect 26712 30598 26740 31622
rect 28920 31580 29296 31589
rect 28976 31578 29000 31580
rect 29056 31578 29080 31580
rect 29136 31578 29160 31580
rect 29216 31578 29240 31580
rect 28976 31526 28986 31578
rect 29230 31526 29240 31578
rect 28976 31524 29000 31526
rect 29056 31524 29080 31526
rect 29136 31524 29160 31526
rect 29216 31524 29240 31526
rect 28920 31515 29296 31524
rect 28180 31036 28556 31045
rect 28236 31034 28260 31036
rect 28316 31034 28340 31036
rect 28396 31034 28420 31036
rect 28476 31034 28500 31036
rect 28236 30982 28246 31034
rect 28490 30982 28500 31034
rect 28236 30980 28260 30982
rect 28316 30980 28340 30982
rect 28396 30980 28420 30982
rect 28476 30980 28500 30982
rect 28180 30971 28556 30980
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 24952 30320 25004 30326
rect 24952 30262 25004 30268
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24780 29850 24808 29990
rect 24768 29844 24820 29850
rect 24768 29786 24820 29792
rect 24964 29714 24992 30262
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 26240 29572 26292 29578
rect 26240 29514 26292 29520
rect 26252 29306 26280 29514
rect 26240 29300 26292 29306
rect 26240 29242 26292 29248
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24032 28960 24084 28966
rect 24032 28902 24084 28908
rect 24044 28082 24072 28902
rect 24032 28076 24084 28082
rect 24032 28018 24084 28024
rect 24032 27872 24084 27878
rect 24032 27814 24084 27820
rect 24044 27713 24072 27814
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 24216 26920 24268 26926
rect 24216 26862 24268 26868
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 24044 26042 24072 26318
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24136 23866 24164 24006
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24124 23656 24176 23662
rect 24124 23598 24176 23604
rect 24136 23186 24164 23598
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 23952 23050 24072 23066
rect 23952 23044 24084 23050
rect 23952 23038 24032 23044
rect 24032 22986 24084 22992
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23952 21146 23980 22578
rect 24044 21962 24072 22986
rect 24124 22568 24176 22574
rect 24228 22556 24256 26862
rect 24320 22964 24348 28970
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24412 26858 24440 26930
rect 24400 26852 24452 26858
rect 24400 26794 24452 26800
rect 24492 26784 24544 26790
rect 24492 26726 24544 26732
rect 24504 25838 24532 26726
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24400 24744 24452 24750
rect 24400 24686 24452 24692
rect 24412 24410 24440 24686
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24412 23118 24440 24346
rect 24504 24290 24532 25774
rect 24688 24682 24716 28970
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24768 26852 24820 26858
rect 24768 26794 24820 26800
rect 24676 24676 24728 24682
rect 24676 24618 24728 24624
rect 24584 24608 24636 24614
rect 24584 24550 24636 24556
rect 24596 24410 24624 24550
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24504 24262 24624 24290
rect 24688 24274 24716 24618
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24400 22976 24452 22982
rect 24320 22936 24400 22964
rect 24400 22918 24452 22924
rect 24176 22528 24256 22556
rect 24124 22510 24176 22516
rect 24032 21956 24084 21962
rect 24032 21898 24084 21904
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 24044 20942 24072 21422
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 23952 20806 23980 20878
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 24044 20466 24072 20878
rect 24136 20602 24164 22510
rect 24412 22166 24440 22918
rect 24504 22778 24532 23258
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 24308 21956 24360 21962
rect 24308 21898 24360 21904
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24228 21350 24256 21490
rect 24320 21350 24348 21898
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24320 21078 24348 21286
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 24412 20942 24440 21286
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24044 19854 24072 20402
rect 24412 20398 24440 20878
rect 24400 20392 24452 20398
rect 24400 20334 24452 20340
rect 24412 19990 24440 20334
rect 24400 19984 24452 19990
rect 24492 19984 24544 19990
rect 24400 19926 24452 19932
rect 24490 19952 24492 19961
rect 24544 19952 24546 19961
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 24412 19174 24440 19926
rect 24490 19887 24546 19896
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18358 24440 19110
rect 24504 18970 24532 19790
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24400 18352 24452 18358
rect 24400 18294 24452 18300
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 23768 17326 23888 17354
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23572 16720 23624 16726
rect 23572 16662 23624 16668
rect 23584 16250 23612 16662
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23480 12776 23532 12782
rect 23480 12718 23532 12724
rect 23388 12232 23440 12238
rect 23202 12200 23258 12209
rect 23112 12164 23164 12170
rect 23388 12174 23440 12180
rect 23202 12135 23258 12144
rect 23112 12106 23164 12112
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 22920 11996 23296 12005
rect 22976 11994 23000 11996
rect 23056 11994 23080 11996
rect 23136 11994 23160 11996
rect 23216 11994 23240 11996
rect 22976 11942 22986 11994
rect 23230 11942 23240 11994
rect 22976 11940 23000 11942
rect 23056 11940 23080 11942
rect 23136 11940 23160 11942
rect 23216 11940 23240 11942
rect 22920 11931 23296 11940
rect 23400 11762 23428 12038
rect 23492 11898 23520 12718
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12442 23704 12582
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23584 12102 23612 12378
rect 23572 12096 23624 12102
rect 23624 12044 23704 12050
rect 23572 12038 23704 12044
rect 23584 12022 23704 12038
rect 23570 11928 23626 11937
rect 23480 11892 23532 11898
rect 23570 11863 23626 11872
rect 23480 11834 23532 11840
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 22920 10908 23296 10917
rect 22976 10906 23000 10908
rect 23056 10906 23080 10908
rect 23136 10906 23160 10908
rect 23216 10906 23240 10908
rect 22976 10854 22986 10906
rect 23230 10854 23240 10906
rect 22976 10852 23000 10854
rect 23056 10852 23080 10854
rect 23136 10852 23160 10854
rect 23216 10852 23240 10854
rect 22920 10843 23296 10852
rect 22848 10764 23060 10792
rect 23032 10033 23060 10764
rect 23584 10266 23612 11863
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23018 10024 23074 10033
rect 22744 9988 22796 9994
rect 22796 9948 22876 9976
rect 23018 9959 23074 9968
rect 23572 9988 23624 9994
rect 22744 9930 22796 9936
rect 22742 9688 22798 9697
rect 22742 9623 22798 9632
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22180 9276 22556 9285
rect 22236 9274 22260 9276
rect 22316 9274 22340 9276
rect 22396 9274 22420 9276
rect 22476 9274 22500 9276
rect 22236 9222 22246 9274
rect 22490 9222 22500 9274
rect 22236 9220 22260 9222
rect 22316 9220 22340 9222
rect 22396 9220 22420 9222
rect 22476 9220 22500 9222
rect 22180 9211 22556 9220
rect 22112 8906 22232 8922
rect 22112 8900 22244 8906
rect 22112 8894 22192 8900
rect 22192 8842 22244 8848
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22112 8430 22140 8774
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21652 6798 21680 7686
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20444 6180 20496 6186
rect 20444 6122 20496 6128
rect 20456 5846 20484 6122
rect 20444 5840 20496 5846
rect 20444 5782 20496 5788
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 21008 5710 21036 6598
rect 21560 6458 21588 6598
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 22020 6254 22048 6598
rect 22112 6390 22140 8366
rect 22180 8188 22556 8197
rect 22236 8186 22260 8188
rect 22316 8186 22340 8188
rect 22396 8186 22420 8188
rect 22476 8186 22500 8188
rect 22236 8134 22246 8186
rect 22490 8134 22500 8186
rect 22236 8132 22260 8134
rect 22316 8132 22340 8134
rect 22396 8132 22420 8134
rect 22476 8132 22500 8134
rect 22180 8123 22556 8132
rect 22180 7100 22556 7109
rect 22236 7098 22260 7100
rect 22316 7098 22340 7100
rect 22396 7098 22420 7100
rect 22476 7098 22500 7100
rect 22236 7046 22246 7098
rect 22490 7046 22500 7098
rect 22236 7044 22260 7046
rect 22316 7044 22340 7046
rect 22396 7044 22420 7046
rect 22476 7044 22500 7046
rect 22180 7035 22556 7044
rect 22664 7002 22692 9454
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22652 6792 22704 6798
rect 22756 6780 22784 9623
rect 22704 6752 22784 6780
rect 22652 6734 22704 6740
rect 22468 6724 22520 6730
rect 22468 6666 22520 6672
rect 22480 6458 22508 6666
rect 22652 6656 22704 6662
rect 22848 6644 22876 9948
rect 23572 9930 23624 9936
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 22920 9820 23296 9829
rect 22976 9818 23000 9820
rect 23056 9818 23080 9820
rect 23136 9818 23160 9820
rect 23216 9818 23240 9820
rect 22976 9766 22986 9818
rect 23230 9766 23240 9818
rect 22976 9764 23000 9766
rect 23056 9764 23080 9766
rect 23136 9764 23160 9766
rect 23216 9764 23240 9766
rect 22920 9755 23296 9764
rect 23388 9716 23440 9722
rect 23294 9688 23350 9697
rect 23388 9658 23440 9664
rect 23294 9623 23350 9632
rect 23308 8945 23336 9623
rect 23400 9586 23428 9658
rect 23492 9586 23520 9862
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23400 9178 23428 9522
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23388 8968 23440 8974
rect 23294 8936 23350 8945
rect 23388 8910 23440 8916
rect 23294 8871 23350 8880
rect 22920 8732 23296 8741
rect 22976 8730 23000 8732
rect 23056 8730 23080 8732
rect 23136 8730 23160 8732
rect 23216 8730 23240 8732
rect 22976 8678 22986 8730
rect 23230 8678 23240 8730
rect 22976 8676 23000 8678
rect 23056 8676 23080 8678
rect 23136 8676 23160 8678
rect 23216 8676 23240 8678
rect 22920 8667 23296 8676
rect 22920 7644 23296 7653
rect 22976 7642 23000 7644
rect 23056 7642 23080 7644
rect 23136 7642 23160 7644
rect 23216 7642 23240 7644
rect 22976 7590 22986 7642
rect 23230 7590 23240 7642
rect 22976 7588 23000 7590
rect 23056 7588 23080 7590
rect 23136 7588 23160 7590
rect 23216 7588 23240 7590
rect 22920 7579 23296 7588
rect 22704 6616 22876 6644
rect 22652 6598 22704 6604
rect 22920 6556 23296 6565
rect 22976 6554 23000 6556
rect 23056 6554 23080 6556
rect 23136 6554 23160 6556
rect 23216 6554 23240 6556
rect 22976 6502 22986 6554
rect 23230 6502 23240 6554
rect 22976 6500 23000 6502
rect 23056 6500 23080 6502
rect 23136 6500 23160 6502
rect 23216 6500 23240 6502
rect 22920 6491 23296 6500
rect 22468 6452 22520 6458
rect 22468 6394 22520 6400
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 22008 6248 22060 6254
rect 22008 6190 22060 6196
rect 22020 5914 22048 6190
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22112 5710 22140 6326
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22180 6012 22556 6021
rect 22236 6010 22260 6012
rect 22316 6010 22340 6012
rect 22396 6010 22420 6012
rect 22476 6010 22500 6012
rect 22236 5958 22246 6010
rect 22490 5958 22500 6010
rect 22236 5956 22260 5958
rect 22316 5956 22340 5958
rect 22396 5956 22420 5958
rect 22476 5956 22500 5958
rect 22180 5947 22556 5956
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22204 5370 22232 5510
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 5098 22324 5578
rect 22664 5370 22692 6054
rect 23216 5914 23244 6258
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23400 5794 23428 8910
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8634 23520 8774
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23584 8430 23612 9930
rect 23676 9654 23704 12022
rect 23768 9722 23796 17326
rect 23952 17252 23980 18226
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17338 24072 18022
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 23860 17224 23980 17252
rect 23860 16114 23888 17224
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23952 16794 23980 17070
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 24044 16590 24072 17274
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24308 16516 24360 16522
rect 24308 16458 24360 16464
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23860 15706 23888 16050
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 23848 15020 23900 15026
rect 23848 14962 23900 14968
rect 23860 10674 23888 14962
rect 24136 13938 24164 15370
rect 24320 14958 24348 16458
rect 24412 16114 24440 16594
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24398 15192 24454 15201
rect 24398 15127 24454 15136
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24228 12442 24256 13806
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24044 12152 24072 12378
rect 24320 12238 24348 14894
rect 24412 13938 24440 15127
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24412 12986 24440 13126
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24216 12164 24268 12170
rect 24044 12124 24216 12152
rect 24216 12106 24268 12112
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 24216 9920 24268 9926
rect 24216 9862 24268 9868
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23664 9648 23716 9654
rect 23664 9590 23716 9596
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 9110 24072 9522
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24136 9178 24164 9386
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8498 24072 8774
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 24228 6458 24256 9862
rect 24320 9450 24348 12174
rect 24504 11898 24532 12174
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 9722 24532 10542
rect 24596 9926 24624 24262
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24780 22642 24808 26794
rect 24872 25838 24900 27474
rect 24964 27470 24992 29038
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 27130 26188 27406
rect 26712 27402 26740 30534
rect 28920 30492 29296 30501
rect 28976 30490 29000 30492
rect 29056 30490 29080 30492
rect 29136 30490 29160 30492
rect 29216 30490 29240 30492
rect 28976 30438 28986 30490
rect 29230 30438 29240 30490
rect 28976 30436 29000 30438
rect 29056 30436 29080 30438
rect 29136 30436 29160 30438
rect 29216 30436 29240 30438
rect 28920 30427 29296 30436
rect 28180 29948 28556 29957
rect 28236 29946 28260 29948
rect 28316 29946 28340 29948
rect 28396 29946 28420 29948
rect 28476 29946 28500 29948
rect 28236 29894 28246 29946
rect 28490 29894 28500 29946
rect 28236 29892 28260 29894
rect 28316 29892 28340 29894
rect 28396 29892 28420 29894
rect 28476 29892 28500 29894
rect 28180 29883 28556 29892
rect 28920 29404 29296 29413
rect 28976 29402 29000 29404
rect 29056 29402 29080 29404
rect 29136 29402 29160 29404
rect 29216 29402 29240 29404
rect 28976 29350 28986 29402
rect 29230 29350 29240 29402
rect 28976 29348 29000 29350
rect 29056 29348 29080 29350
rect 29136 29348 29160 29350
rect 29216 29348 29240 29350
rect 28920 29339 29296 29348
rect 28180 28860 28556 28869
rect 28236 28858 28260 28860
rect 28316 28858 28340 28860
rect 28396 28858 28420 28860
rect 28476 28858 28500 28860
rect 28236 28806 28246 28858
rect 28490 28806 28500 28858
rect 28236 28804 28260 28806
rect 28316 28804 28340 28806
rect 28396 28804 28420 28806
rect 28476 28804 28500 28806
rect 28180 28795 28556 28804
rect 28920 28316 29296 28325
rect 28976 28314 29000 28316
rect 29056 28314 29080 28316
rect 29136 28314 29160 28316
rect 29216 28314 29240 28316
rect 28976 28262 28986 28314
rect 29230 28262 29240 28314
rect 28976 28260 29000 28262
rect 29056 28260 29080 28262
rect 29136 28260 29160 28262
rect 29216 28260 29240 28262
rect 28920 28251 29296 28260
rect 28180 27772 28556 27781
rect 28236 27770 28260 27772
rect 28316 27770 28340 27772
rect 28396 27770 28420 27772
rect 28476 27770 28500 27772
rect 28236 27718 28246 27770
rect 28490 27718 28500 27770
rect 28236 27716 28260 27718
rect 28316 27716 28340 27718
rect 28396 27716 28420 27718
rect 28476 27716 28500 27718
rect 28180 27707 28556 27716
rect 26700 27396 26752 27402
rect 26700 27338 26752 27344
rect 27344 27396 27396 27402
rect 27344 27338 27396 27344
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 26344 27130 26372 27270
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 25780 27056 25832 27062
rect 25780 26998 25832 27004
rect 25044 26920 25096 26926
rect 25044 26862 25096 26868
rect 25056 26586 25084 26862
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25792 26518 25820 26998
rect 25780 26512 25832 26518
rect 25780 26454 25832 26460
rect 25792 25906 25820 26454
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24872 24410 24900 25774
rect 25228 24744 25280 24750
rect 25228 24686 25280 24692
rect 24860 24404 24912 24410
rect 24860 24346 24912 24352
rect 25240 23526 25268 24686
rect 25596 24064 25648 24070
rect 25596 24006 25648 24012
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 25608 23866 25636 24006
rect 25976 23866 26004 24006
rect 25596 23860 25648 23866
rect 25596 23802 25648 23808
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 26332 23656 26384 23662
rect 26332 23598 26384 23604
rect 25228 23520 25280 23526
rect 25228 23462 25280 23468
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24688 18902 24716 20402
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18086 24716 18566
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24780 17678 24808 19654
rect 25056 19378 25084 23054
rect 25240 23050 25268 23462
rect 26344 23322 26372 23598
rect 26516 23520 26568 23526
rect 26516 23462 26568 23468
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26528 23118 26556 23462
rect 26516 23112 26568 23118
rect 26516 23054 26568 23060
rect 25228 23044 25280 23050
rect 25228 22986 25280 22992
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 26620 19446 26648 19654
rect 26608 19440 26660 19446
rect 26608 19382 26660 19388
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24872 18154 24900 18566
rect 24964 18290 24992 19314
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24860 18148 24912 18154
rect 24860 18090 24912 18096
rect 25056 17746 25084 19314
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25332 18970 25360 19246
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25136 18760 25188 18766
rect 25136 18702 25188 18708
rect 25148 17882 25176 18702
rect 26712 18222 26740 19790
rect 26700 18216 26752 18222
rect 26700 18158 26752 18164
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 26344 17882 26372 18022
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 24780 17338 24808 17614
rect 25516 17338 25544 17614
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25504 17332 25556 17338
rect 25504 17274 25556 17280
rect 24780 16590 24808 17274
rect 24860 17060 24912 17066
rect 24860 17002 24912 17008
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24872 16250 24900 17002
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 25516 16794 25544 16934
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24688 13394 24716 14758
rect 25516 14074 25544 16118
rect 26148 16108 26200 16114
rect 26148 16050 26200 16056
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25700 15026 25728 15846
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25884 14822 25912 15506
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26068 14958 26096 15438
rect 26160 15162 26188 16050
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 26068 14618 26096 14894
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24492 9716 24544 9722
rect 24492 9658 24544 9664
rect 24688 9602 24716 13330
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12918 24808 13126
rect 25792 12986 25820 13262
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 24768 12912 24820 12918
rect 24768 12854 24820 12860
rect 25240 12102 25268 12922
rect 25884 12782 25912 13466
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25780 11076 25832 11082
rect 25780 11018 25832 11024
rect 25792 10810 25820 11018
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9722 24900 9862
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24412 9574 24716 9602
rect 24768 9580 24820 9586
rect 24412 9518 24440 9574
rect 24768 9522 24820 9528
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 24308 6724 24360 6730
rect 24308 6666 24360 6672
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 22848 5766 23428 5794
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 22848 5166 22876 5766
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 22920 5468 23296 5477
rect 22976 5466 23000 5468
rect 23056 5466 23080 5468
rect 23136 5466 23160 5468
rect 23216 5466 23240 5468
rect 22976 5414 22986 5466
rect 23230 5414 23240 5466
rect 22976 5412 23000 5414
rect 23056 5412 23080 5414
rect 23136 5412 23160 5414
rect 23216 5412 23240 5414
rect 22920 5403 23296 5412
rect 23400 5370 23428 5578
rect 23584 5574 23612 6394
rect 24320 6186 24348 6666
rect 24412 6322 24440 9454
rect 24780 9110 24808 9522
rect 24964 9450 24992 10066
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24596 6798 24624 9046
rect 24872 6798 24900 9386
rect 24964 8634 24992 9386
rect 25056 9178 25084 9998
rect 25412 9920 25464 9926
rect 25412 9862 25464 9868
rect 25424 9722 25452 9862
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25884 9518 25912 12718
rect 26160 12170 26188 14962
rect 26252 14414 26280 16594
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26528 16114 26556 16390
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26712 15706 26740 15846
rect 26700 15700 26752 15706
rect 26700 15642 26752 15648
rect 26516 15496 26568 15502
rect 26516 15438 26568 15444
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26344 14482 26372 14894
rect 26332 14476 26384 14482
rect 26332 14418 26384 14424
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26252 12306 26280 14350
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26148 12164 26200 12170
rect 26148 12106 26200 12112
rect 26344 11558 26372 14418
rect 26436 12986 26464 14962
rect 26528 14890 26556 15438
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26712 15162 26740 15302
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26516 14884 26568 14890
rect 26516 14826 26568 14832
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26700 12776 26752 12782
rect 26700 12718 26752 12724
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26436 12238 26464 12582
rect 26712 12442 26740 12718
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26804 12322 26832 14758
rect 26620 12294 26832 12322
rect 26620 12238 26648 12294
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26700 12232 26752 12238
rect 26896 12186 26924 24006
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17202 27016 18158
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 27080 17610 27108 18022
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26988 15434 27016 17138
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 27172 16590 27200 16934
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 26700 12174 26752 12180
rect 26436 11898 26464 12174
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 26436 11354 26464 11698
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26424 11348 26476 11354
rect 26424 11290 26476 11296
rect 26436 9518 26464 11290
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25872 9512 25924 9518
rect 25872 9454 25924 9460
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 25044 9172 25096 9178
rect 25044 9114 25096 9120
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25148 6798 25176 8871
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24860 6792 24912 6798
rect 24860 6734 24912 6740
rect 25136 6792 25188 6798
rect 25136 6734 25188 6740
rect 24768 6724 24820 6730
rect 24768 6666 24820 6672
rect 24780 6458 24808 6666
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24308 6180 24360 6186
rect 24308 6122 24360 6128
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24216 6112 24268 6118
rect 24216 6054 24268 6060
rect 24136 5914 24164 6054
rect 24228 5914 24256 6054
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 23676 5302 23704 5510
rect 24320 5370 24348 6122
rect 24688 5658 24716 6394
rect 24780 5914 24808 6394
rect 25424 6186 25452 9454
rect 25596 9376 25648 9382
rect 25596 9318 25648 9324
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 25608 9178 25636 9318
rect 26068 9178 26096 9318
rect 25596 9172 25648 9178
rect 25596 9114 25648 9120
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25792 8634 25820 8774
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25884 8498 25912 8774
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 25412 5840 25464 5846
rect 25412 5782 25464 5788
rect 24688 5642 24808 5658
rect 24688 5636 24820 5642
rect 24688 5630 24768 5636
rect 24768 5578 24820 5584
rect 24308 5364 24360 5370
rect 24308 5306 24360 5312
rect 23664 5296 23716 5302
rect 25424 5250 25452 5782
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 23664 5238 23716 5244
rect 25332 5234 25452 5250
rect 25516 5234 25544 5646
rect 25320 5228 25452 5234
rect 25372 5222 25452 5228
rect 25504 5228 25556 5234
rect 25320 5170 25372 5176
rect 25504 5170 25556 5176
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 22284 5092 22336 5098
rect 22284 5034 22336 5040
rect 22180 4924 22556 4933
rect 22236 4922 22260 4924
rect 22316 4922 22340 4924
rect 22396 4922 22420 4924
rect 22476 4922 22500 4924
rect 22236 4870 22246 4922
rect 22490 4870 22500 4922
rect 22236 4868 22260 4870
rect 22316 4868 22340 4870
rect 22396 4868 22420 4870
rect 22476 4868 22500 4870
rect 22180 4859 22556 4868
rect 22920 4380 23296 4389
rect 22976 4378 23000 4380
rect 23056 4378 23080 4380
rect 23136 4378 23160 4380
rect 23216 4378 23240 4380
rect 22976 4326 22986 4378
rect 23230 4326 23240 4378
rect 22976 4324 23000 4326
rect 23056 4324 23080 4326
rect 23136 4324 23160 4326
rect 23216 4324 23240 4326
rect 22920 4315 23296 4324
rect 25516 4146 25544 5170
rect 26252 4622 26280 6598
rect 26528 5778 26556 11494
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26620 5030 26648 12174
rect 26712 5234 26740 12174
rect 26804 12158 26924 12186
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 26804 11354 26832 12158
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26896 11354 26924 12038
rect 26988 11694 27016 12174
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 26792 11348 26844 11354
rect 26792 11290 26844 11296
rect 26884 11348 26936 11354
rect 26884 11290 26936 11296
rect 27080 11132 27108 16050
rect 27264 15162 27292 27270
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27172 14414 27200 14894
rect 27252 14816 27304 14822
rect 27252 14758 27304 14764
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27264 14346 27292 14758
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27356 11150 27384 27338
rect 28920 27228 29296 27237
rect 28976 27226 29000 27228
rect 29056 27226 29080 27228
rect 29136 27226 29160 27228
rect 29216 27226 29240 27228
rect 28976 27174 28986 27226
rect 29230 27174 29240 27226
rect 28976 27172 29000 27174
rect 29056 27172 29080 27174
rect 29136 27172 29160 27174
rect 29216 27172 29240 27174
rect 28920 27163 29296 27172
rect 28180 26684 28556 26693
rect 28236 26682 28260 26684
rect 28316 26682 28340 26684
rect 28396 26682 28420 26684
rect 28476 26682 28500 26684
rect 28236 26630 28246 26682
rect 28490 26630 28500 26682
rect 28236 26628 28260 26630
rect 28316 26628 28340 26630
rect 28396 26628 28420 26630
rect 28476 26628 28500 26630
rect 28180 26619 28556 26628
rect 28920 26140 29296 26149
rect 28976 26138 29000 26140
rect 29056 26138 29080 26140
rect 29136 26138 29160 26140
rect 29216 26138 29240 26140
rect 28976 26086 28986 26138
rect 29230 26086 29240 26138
rect 28976 26084 29000 26086
rect 29056 26084 29080 26086
rect 29136 26084 29160 26086
rect 29216 26084 29240 26086
rect 28920 26075 29296 26084
rect 28180 25596 28556 25605
rect 28236 25594 28260 25596
rect 28316 25594 28340 25596
rect 28396 25594 28420 25596
rect 28476 25594 28500 25596
rect 28236 25542 28246 25594
rect 28490 25542 28500 25594
rect 28236 25540 28260 25542
rect 28316 25540 28340 25542
rect 28396 25540 28420 25542
rect 28476 25540 28500 25542
rect 28180 25531 28556 25540
rect 31300 25424 31352 25430
rect 31300 25366 31352 25372
rect 30656 25288 30708 25294
rect 31312 25265 31340 25366
rect 30656 25230 30708 25236
rect 31298 25256 31354 25265
rect 28920 25052 29296 25061
rect 28976 25050 29000 25052
rect 29056 25050 29080 25052
rect 29136 25050 29160 25052
rect 29216 25050 29240 25052
rect 28976 24998 28986 25050
rect 29230 24998 29240 25050
rect 28976 24996 29000 24998
rect 29056 24996 29080 24998
rect 29136 24996 29160 24998
rect 29216 24996 29240 24998
rect 28920 24987 29296 24996
rect 28180 24508 28556 24517
rect 28236 24506 28260 24508
rect 28316 24506 28340 24508
rect 28396 24506 28420 24508
rect 28476 24506 28500 24508
rect 28236 24454 28246 24506
rect 28490 24454 28500 24506
rect 28236 24452 28260 24454
rect 28316 24452 28340 24454
rect 28396 24452 28420 24454
rect 28476 24452 28500 24454
rect 28180 24443 28556 24452
rect 28920 23964 29296 23973
rect 28976 23962 29000 23964
rect 29056 23962 29080 23964
rect 29136 23962 29160 23964
rect 29216 23962 29240 23964
rect 28976 23910 28986 23962
rect 29230 23910 29240 23962
rect 28976 23908 29000 23910
rect 29056 23908 29080 23910
rect 29136 23908 29160 23910
rect 29216 23908 29240 23910
rect 28920 23899 29296 23908
rect 28180 23420 28556 23429
rect 28236 23418 28260 23420
rect 28316 23418 28340 23420
rect 28396 23418 28420 23420
rect 28476 23418 28500 23420
rect 28236 23366 28246 23418
rect 28490 23366 28500 23418
rect 28236 23364 28260 23366
rect 28316 23364 28340 23366
rect 28396 23364 28420 23366
rect 28476 23364 28500 23366
rect 28180 23355 28556 23364
rect 28920 22876 29296 22885
rect 28976 22874 29000 22876
rect 29056 22874 29080 22876
rect 29136 22874 29160 22876
rect 29216 22874 29240 22876
rect 28976 22822 28986 22874
rect 29230 22822 29240 22874
rect 28976 22820 29000 22822
rect 29056 22820 29080 22822
rect 29136 22820 29160 22822
rect 29216 22820 29240 22822
rect 28920 22811 29296 22820
rect 28180 22332 28556 22341
rect 28236 22330 28260 22332
rect 28316 22330 28340 22332
rect 28396 22330 28420 22332
rect 28476 22330 28500 22332
rect 28236 22278 28246 22330
rect 28490 22278 28500 22330
rect 28236 22276 28260 22278
rect 28316 22276 28340 22278
rect 28396 22276 28420 22278
rect 28476 22276 28500 22278
rect 28180 22267 28556 22276
rect 28920 21788 29296 21797
rect 28976 21786 29000 21788
rect 29056 21786 29080 21788
rect 29136 21786 29160 21788
rect 29216 21786 29240 21788
rect 28976 21734 28986 21786
rect 29230 21734 29240 21786
rect 28976 21732 29000 21734
rect 29056 21732 29080 21734
rect 29136 21732 29160 21734
rect 29216 21732 29240 21734
rect 28920 21723 29296 21732
rect 28180 21244 28556 21253
rect 28236 21242 28260 21244
rect 28316 21242 28340 21244
rect 28396 21242 28420 21244
rect 28476 21242 28500 21244
rect 28236 21190 28246 21242
rect 28490 21190 28500 21242
rect 28236 21188 28260 21190
rect 28316 21188 28340 21190
rect 28396 21188 28420 21190
rect 28476 21188 28500 21190
rect 28180 21179 28556 21188
rect 28920 20700 29296 20709
rect 28976 20698 29000 20700
rect 29056 20698 29080 20700
rect 29136 20698 29160 20700
rect 29216 20698 29240 20700
rect 28976 20646 28986 20698
rect 29230 20646 29240 20698
rect 28976 20644 29000 20646
rect 29056 20644 29080 20646
rect 29136 20644 29160 20646
rect 29216 20644 29240 20646
rect 28920 20635 29296 20644
rect 28180 20156 28556 20165
rect 28236 20154 28260 20156
rect 28316 20154 28340 20156
rect 28396 20154 28420 20156
rect 28476 20154 28500 20156
rect 28236 20102 28246 20154
rect 28490 20102 28500 20154
rect 28236 20100 28260 20102
rect 28316 20100 28340 20102
rect 28396 20100 28420 20102
rect 28476 20100 28500 20102
rect 28180 20091 28556 20100
rect 28920 19612 29296 19621
rect 28976 19610 29000 19612
rect 29056 19610 29080 19612
rect 29136 19610 29160 19612
rect 29216 19610 29240 19612
rect 28976 19558 28986 19610
rect 29230 19558 29240 19610
rect 28976 19556 29000 19558
rect 29056 19556 29080 19558
rect 29136 19556 29160 19558
rect 29216 19556 29240 19558
rect 28920 19547 29296 19556
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 28180 19068 28556 19077
rect 28236 19066 28260 19068
rect 28316 19066 28340 19068
rect 28396 19066 28420 19068
rect 28476 19066 28500 19068
rect 28236 19014 28246 19066
rect 28490 19014 28500 19066
rect 28236 19012 28260 19014
rect 28316 19012 28340 19014
rect 28396 19012 28420 19014
rect 28476 19012 28500 19014
rect 28180 19003 28556 19012
rect 28920 18524 29296 18533
rect 28976 18522 29000 18524
rect 29056 18522 29080 18524
rect 29136 18522 29160 18524
rect 29216 18522 29240 18524
rect 28976 18470 28986 18522
rect 29230 18470 29240 18522
rect 28976 18468 29000 18470
rect 29056 18468 29080 18470
rect 29136 18468 29160 18470
rect 29216 18468 29240 18470
rect 28920 18459 29296 18468
rect 27620 18080 27672 18086
rect 27620 18022 27672 18028
rect 27632 16794 27660 18022
rect 28180 17980 28556 17989
rect 28236 17978 28260 17980
rect 28316 17978 28340 17980
rect 28396 17978 28420 17980
rect 28476 17978 28500 17980
rect 28236 17926 28246 17978
rect 28490 17926 28500 17978
rect 28236 17924 28260 17926
rect 28316 17924 28340 17926
rect 28396 17924 28420 17926
rect 28476 17924 28500 17926
rect 28180 17915 28556 17924
rect 28920 17436 29296 17445
rect 28976 17434 29000 17436
rect 29056 17434 29080 17436
rect 29136 17434 29160 17436
rect 29216 17434 29240 17436
rect 28976 17382 28986 17434
rect 29230 17382 29240 17434
rect 28976 17380 29000 17382
rect 29056 17380 29080 17382
rect 29136 17380 29160 17382
rect 29216 17380 29240 17382
rect 28920 17371 29296 17380
rect 28180 16892 28556 16901
rect 28236 16890 28260 16892
rect 28316 16890 28340 16892
rect 28396 16890 28420 16892
rect 28476 16890 28500 16892
rect 28236 16838 28246 16890
rect 28490 16838 28500 16890
rect 28236 16836 28260 16838
rect 28316 16836 28340 16838
rect 28396 16836 28420 16838
rect 28476 16836 28500 16838
rect 28180 16827 28556 16836
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 28920 16348 29296 16357
rect 28976 16346 29000 16348
rect 29056 16346 29080 16348
rect 29136 16346 29160 16348
rect 29216 16346 29240 16348
rect 28976 16294 28986 16346
rect 29230 16294 29240 16346
rect 28976 16292 29000 16294
rect 29056 16292 29080 16294
rect 29136 16292 29160 16294
rect 29216 16292 29240 16294
rect 28920 16283 29296 16292
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27540 15706 27568 15982
rect 28180 15804 28556 15813
rect 28236 15802 28260 15804
rect 28316 15802 28340 15804
rect 28396 15802 28420 15804
rect 28476 15802 28500 15804
rect 28236 15750 28246 15802
rect 28490 15750 28500 15802
rect 28236 15748 28260 15750
rect 28316 15748 28340 15750
rect 28396 15748 28420 15750
rect 28476 15748 28500 15750
rect 28180 15739 28556 15748
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 29656 15570 29684 19314
rect 29644 15564 29696 15570
rect 29644 15506 29696 15512
rect 27436 15428 27488 15434
rect 27436 15370 27488 15376
rect 27160 11144 27212 11150
rect 27080 11104 27160 11132
rect 27160 11086 27212 11092
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 27068 5704 27120 5710
rect 27068 5646 27120 5652
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 27080 5166 27108 5646
rect 27068 5160 27120 5166
rect 27068 5102 27120 5108
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 27172 4622 27200 11086
rect 27448 5114 27476 15370
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27816 15094 27844 15302
rect 28920 15260 29296 15269
rect 28976 15258 29000 15260
rect 29056 15258 29080 15260
rect 29136 15258 29160 15260
rect 29216 15258 29240 15260
rect 28976 15206 28986 15258
rect 29230 15206 29240 15258
rect 28976 15204 29000 15206
rect 29056 15204 29080 15206
rect 29136 15204 29160 15206
rect 29216 15204 29240 15206
rect 28920 15195 29296 15204
rect 29656 15162 29684 15506
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 29368 14952 29420 14958
rect 29368 14894 29420 14900
rect 28180 14716 28556 14725
rect 28236 14714 28260 14716
rect 28316 14714 28340 14716
rect 28396 14714 28420 14716
rect 28476 14714 28500 14716
rect 28236 14662 28246 14714
rect 28490 14662 28500 14714
rect 28236 14660 28260 14662
rect 28316 14660 28340 14662
rect 28396 14660 28420 14662
rect 28476 14660 28500 14662
rect 28180 14651 28556 14660
rect 28920 14172 29296 14181
rect 28976 14170 29000 14172
rect 29056 14170 29080 14172
rect 29136 14170 29160 14172
rect 29216 14170 29240 14172
rect 28976 14118 28986 14170
rect 29230 14118 29240 14170
rect 28976 14116 29000 14118
rect 29056 14116 29080 14118
rect 29136 14116 29160 14118
rect 29216 14116 29240 14118
rect 28920 14107 29296 14116
rect 28180 13628 28556 13637
rect 28236 13626 28260 13628
rect 28316 13626 28340 13628
rect 28396 13626 28420 13628
rect 28476 13626 28500 13628
rect 28236 13574 28246 13626
rect 28490 13574 28500 13626
rect 28236 13572 28260 13574
rect 28316 13572 28340 13574
rect 28396 13572 28420 13574
rect 28476 13572 28500 13574
rect 28180 13563 28556 13572
rect 29380 13530 29408 14894
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 28920 13084 29296 13093
rect 28976 13082 29000 13084
rect 29056 13082 29080 13084
rect 29136 13082 29160 13084
rect 29216 13082 29240 13084
rect 28976 13030 28986 13082
rect 29230 13030 29240 13082
rect 28976 13028 29000 13030
rect 29056 13028 29080 13030
rect 29136 13028 29160 13030
rect 29216 13028 29240 13030
rect 28920 13019 29296 13028
rect 29380 12986 29408 13466
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27632 11354 27660 12106
rect 28092 11898 28120 12718
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28180 12540 28556 12549
rect 28236 12538 28260 12540
rect 28316 12538 28340 12540
rect 28396 12538 28420 12540
rect 28476 12538 28500 12540
rect 28236 12486 28246 12538
rect 28490 12486 28500 12538
rect 28236 12484 28260 12486
rect 28316 12484 28340 12486
rect 28396 12484 28420 12486
rect 28476 12484 28500 12486
rect 28180 12475 28556 12484
rect 28644 12170 28672 12582
rect 30668 12442 30696 25230
rect 31298 25191 31354 25200
rect 30932 19168 30984 19174
rect 30930 19136 30932 19145
rect 30984 19136 30986 19145
rect 30930 19071 30986 19080
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31312 13025 31340 13194
rect 31298 13016 31354 13025
rect 31298 12951 31354 12960
rect 30656 12436 30708 12442
rect 30656 12378 30708 12384
rect 28632 12164 28684 12170
rect 28632 12106 28684 12112
rect 28920 11996 29296 12005
rect 28976 11994 29000 11996
rect 29056 11994 29080 11996
rect 29136 11994 29160 11996
rect 29216 11994 29240 11996
rect 28976 11942 28986 11994
rect 29230 11942 29240 11994
rect 28976 11940 29000 11942
rect 29056 11940 29080 11942
rect 29136 11940 29160 11942
rect 29216 11940 29240 11942
rect 28920 11931 29296 11940
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 30668 11762 30696 12378
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27724 11354 27752 11494
rect 28180 11452 28556 11461
rect 28236 11450 28260 11452
rect 28316 11450 28340 11452
rect 28396 11450 28420 11452
rect 28476 11450 28500 11452
rect 28236 11398 28246 11450
rect 28490 11398 28500 11450
rect 28236 11396 28260 11398
rect 28316 11396 28340 11398
rect 28396 11396 28420 11398
rect 28476 11396 28500 11398
rect 28180 11387 28556 11396
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 28920 10908 29296 10917
rect 28976 10906 29000 10908
rect 29056 10906 29080 10908
rect 29136 10906 29160 10908
rect 29216 10906 29240 10908
rect 28976 10854 28986 10906
rect 29230 10854 29240 10906
rect 28976 10852 29000 10854
rect 29056 10852 29080 10854
rect 29136 10852 29160 10854
rect 29216 10852 29240 10854
rect 28920 10843 29296 10852
rect 28180 10364 28556 10373
rect 28236 10362 28260 10364
rect 28316 10362 28340 10364
rect 28396 10362 28420 10364
rect 28476 10362 28500 10364
rect 28236 10310 28246 10362
rect 28490 10310 28500 10362
rect 28236 10308 28260 10310
rect 28316 10308 28340 10310
rect 28396 10308 28420 10310
rect 28476 10308 28500 10310
rect 28180 10299 28556 10308
rect 28920 9820 29296 9829
rect 28976 9818 29000 9820
rect 29056 9818 29080 9820
rect 29136 9818 29160 9820
rect 29216 9818 29240 9820
rect 28976 9766 28986 9818
rect 29230 9766 29240 9818
rect 28976 9764 29000 9766
rect 29056 9764 29080 9766
rect 29136 9764 29160 9766
rect 29216 9764 29240 9766
rect 28920 9755 29296 9764
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 28180 9276 28556 9285
rect 28236 9274 28260 9276
rect 28316 9274 28340 9276
rect 28396 9274 28420 9276
rect 28476 9274 28500 9276
rect 28236 9222 28246 9274
rect 28490 9222 28500 9274
rect 28236 9220 28260 9222
rect 28316 9220 28340 9222
rect 28396 9220 28420 9222
rect 28476 9220 28500 9222
rect 28180 9211 28556 9220
rect 28920 8732 29296 8741
rect 28976 8730 29000 8732
rect 29056 8730 29080 8732
rect 29136 8730 29160 8732
rect 29216 8730 29240 8732
rect 28976 8678 28986 8730
rect 29230 8678 29240 8730
rect 28976 8676 29000 8678
rect 29056 8676 29080 8678
rect 29136 8676 29160 8678
rect 29216 8676 29240 8678
rect 28920 8667 29296 8676
rect 28180 8188 28556 8197
rect 28236 8186 28260 8188
rect 28316 8186 28340 8188
rect 28396 8186 28420 8188
rect 28476 8186 28500 8188
rect 28236 8134 28246 8186
rect 28490 8134 28500 8186
rect 28236 8132 28260 8134
rect 28316 8132 28340 8134
rect 28396 8132 28420 8134
rect 28476 8132 28500 8134
rect 28180 8123 28556 8132
rect 30760 8090 30788 9522
rect 30748 8084 30800 8090
rect 30748 8026 30800 8032
rect 31300 7880 31352 7886
rect 31300 7822 31352 7828
rect 28920 7644 29296 7653
rect 28976 7642 29000 7644
rect 29056 7642 29080 7644
rect 29136 7642 29160 7644
rect 29216 7642 29240 7644
rect 28976 7590 28986 7642
rect 29230 7590 29240 7642
rect 28976 7588 29000 7590
rect 29056 7588 29080 7590
rect 29136 7588 29160 7590
rect 29216 7588 29240 7590
rect 28920 7579 29296 7588
rect 31312 7585 31340 7822
rect 31298 7576 31354 7585
rect 31298 7511 31354 7520
rect 28180 7100 28556 7109
rect 28236 7098 28260 7100
rect 28316 7098 28340 7100
rect 28396 7098 28420 7100
rect 28476 7098 28500 7100
rect 28236 7046 28246 7098
rect 28490 7046 28500 7098
rect 28236 7044 28260 7046
rect 28316 7044 28340 7046
rect 28396 7044 28420 7046
rect 28476 7044 28500 7046
rect 28180 7035 28556 7044
rect 28920 6556 29296 6565
rect 28976 6554 29000 6556
rect 29056 6554 29080 6556
rect 29136 6554 29160 6556
rect 29216 6554 29240 6556
rect 28976 6502 28986 6554
rect 29230 6502 29240 6554
rect 28976 6500 29000 6502
rect 29056 6500 29080 6502
rect 29136 6500 29160 6502
rect 29216 6500 29240 6502
rect 28920 6491 29296 6500
rect 28180 6012 28556 6021
rect 28236 6010 28260 6012
rect 28316 6010 28340 6012
rect 28396 6010 28420 6012
rect 28476 6010 28500 6012
rect 28236 5958 28246 6010
rect 28490 5958 28500 6010
rect 28236 5956 28260 5958
rect 28316 5956 28340 5958
rect 28396 5956 28420 5958
rect 28476 5956 28500 5958
rect 28180 5947 28556 5956
rect 28920 5468 29296 5477
rect 28976 5466 29000 5468
rect 29056 5466 29080 5468
rect 29136 5466 29160 5468
rect 29216 5466 29240 5468
rect 28976 5414 28986 5466
rect 29230 5414 29240 5466
rect 28976 5412 29000 5414
rect 29056 5412 29080 5414
rect 29136 5412 29160 5414
rect 29216 5412 29240 5414
rect 28920 5403 29296 5412
rect 27356 5086 27476 5114
rect 26240 4616 26292 4622
rect 26240 4558 26292 4564
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 3398 19472 4014
rect 22180 3836 22556 3845
rect 22236 3834 22260 3836
rect 22316 3834 22340 3836
rect 22396 3834 22420 3836
rect 22476 3834 22500 3836
rect 22236 3782 22246 3834
rect 22490 3782 22500 3834
rect 22236 3780 22260 3782
rect 22316 3780 22340 3782
rect 22396 3780 22420 3782
rect 22476 3780 22500 3782
rect 22180 3771 22556 3780
rect 27356 3670 27384 5086
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27448 4826 27476 4966
rect 28180 4924 28556 4933
rect 28236 4922 28260 4924
rect 28316 4922 28340 4924
rect 28396 4922 28420 4924
rect 28476 4922 28500 4924
rect 28236 4870 28246 4922
rect 28490 4870 28500 4922
rect 28236 4868 28260 4870
rect 28316 4868 28340 4870
rect 28396 4868 28420 4870
rect 28476 4868 28500 4870
rect 28180 4859 28556 4868
rect 27436 4820 27488 4826
rect 27436 4762 27488 4768
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27632 4078 27660 4422
rect 27712 4208 27764 4214
rect 27712 4150 27764 4156
rect 27620 4072 27672 4078
rect 27620 4014 27672 4020
rect 27724 3738 27752 4150
rect 28736 3942 28764 4558
rect 28920 4380 29296 4389
rect 28976 4378 29000 4380
rect 29056 4378 29080 4380
rect 29136 4378 29160 4380
rect 29216 4378 29240 4380
rect 28976 4326 28986 4378
rect 29230 4326 29240 4378
rect 28976 4324 29000 4326
rect 29056 4324 29080 4326
rect 29136 4324 29160 4326
rect 29216 4324 29240 4326
rect 28920 4315 29296 4324
rect 28724 3936 28776 3942
rect 28724 3878 28776 3884
rect 28180 3836 28556 3845
rect 28236 3834 28260 3836
rect 28316 3834 28340 3836
rect 28396 3834 28420 3836
rect 28476 3834 28500 3836
rect 28236 3782 28246 3834
rect 28490 3782 28500 3834
rect 28236 3780 28260 3782
rect 28316 3780 28340 3782
rect 28396 3780 28420 3782
rect 28476 3780 28500 3782
rect 28180 3771 28556 3780
rect 27712 3732 27764 3738
rect 27712 3674 27764 3680
rect 27344 3664 27396 3670
rect 27344 3606 27396 3612
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 16180 2748 16556 2757
rect 16236 2746 16260 2748
rect 16316 2746 16340 2748
rect 16396 2746 16420 2748
rect 16476 2746 16500 2748
rect 18984 2746 19196 2774
rect 16236 2694 16246 2746
rect 16490 2694 16500 2746
rect 16236 2692 16260 2694
rect 16316 2692 16340 2694
rect 16396 2692 16420 2694
rect 16476 2692 16500 2694
rect 16180 2683 16556 2692
rect 19168 2446 19196 2746
rect 20272 2446 20300 3334
rect 22920 3292 23296 3301
rect 22976 3290 23000 3292
rect 23056 3290 23080 3292
rect 23136 3290 23160 3292
rect 23216 3290 23240 3292
rect 22976 3238 22986 3290
rect 23230 3238 23240 3290
rect 22976 3236 23000 3238
rect 23056 3236 23080 3238
rect 23136 3236 23160 3238
rect 23216 3236 23240 3238
rect 22920 3227 23296 3236
rect 22180 2748 22556 2757
rect 22236 2746 22260 2748
rect 22316 2746 22340 2748
rect 22396 2746 22420 2748
rect 22476 2746 22500 2748
rect 22236 2694 22246 2746
rect 22490 2694 22500 2746
rect 22236 2692 22260 2694
rect 22316 2692 22340 2694
rect 22396 2692 22420 2694
rect 22476 2692 22500 2694
rect 22180 2683 22556 2692
rect 28180 2748 28556 2757
rect 28236 2746 28260 2748
rect 28316 2746 28340 2748
rect 28396 2746 28420 2748
rect 28476 2746 28500 2748
rect 28236 2694 28246 2746
rect 28490 2694 28500 2746
rect 28236 2692 28260 2694
rect 28316 2692 28340 2694
rect 28396 2692 28420 2694
rect 28476 2692 28500 2694
rect 28180 2683 28556 2692
rect 28736 2446 28764 3878
rect 28920 3292 29296 3301
rect 28976 3290 29000 3292
rect 29056 3290 29080 3292
rect 29136 3290 29160 3292
rect 29216 3290 29240 3292
rect 28976 3238 28986 3290
rect 29230 3238 29240 3290
rect 28976 3236 29000 3238
rect 29056 3236 29080 3238
rect 29136 3236 29160 3238
rect 29216 3236 29240 3238
rect 28920 3227 29296 3236
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 10796 2372 10928 2378
rect 10796 2366 10876 2372
rect 32 800 60 2314
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 4920 2204 5296 2213
rect 4976 2202 5000 2204
rect 5056 2202 5080 2204
rect 5136 2202 5160 2204
rect 5216 2202 5240 2204
rect 4976 2150 4986 2202
rect 5230 2150 5240 2202
rect 4976 2148 5000 2150
rect 5056 2148 5080 2150
rect 5136 2148 5160 2150
rect 5216 2148 5240 2150
rect 4920 2139 5296 2148
rect 5368 1170 5396 2246
rect 5184 1142 5396 1170
rect 10796 1170 10824 2366
rect 10876 2314 10928 2320
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 28540 2372 28592 2378
rect 28540 2314 28592 2320
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 10920 2204 11296 2213
rect 10976 2202 11000 2204
rect 11056 2202 11080 2204
rect 11136 2202 11160 2204
rect 11216 2202 11240 2204
rect 10976 2150 10986 2202
rect 11230 2150 11240 2202
rect 10976 2148 11000 2150
rect 11056 2148 11080 2150
rect 11136 2148 11160 2150
rect 11216 2148 11240 2150
rect 10920 2139 11296 2148
rect 10796 1142 11008 1170
rect 5184 800 5212 1142
rect 10980 800 11008 1142
rect 16776 800 16804 2246
rect 16920 2204 17296 2213
rect 16976 2202 17000 2204
rect 17056 2202 17080 2204
rect 17136 2202 17160 2204
rect 17216 2202 17240 2204
rect 16976 2150 16986 2202
rect 17230 2150 17240 2202
rect 16976 2148 17000 2150
rect 17056 2148 17080 2150
rect 17136 2148 17160 2150
rect 17216 2148 17240 2150
rect 16920 2139 17296 2148
rect 22572 800 22600 2246
rect 22920 2204 23296 2213
rect 22976 2202 23000 2204
rect 23056 2202 23080 2204
rect 23136 2202 23160 2204
rect 23216 2202 23240 2204
rect 22976 2150 22986 2202
rect 23230 2150 23240 2202
rect 22976 2148 23000 2150
rect 23056 2148 23080 2150
rect 23136 2148 23160 2150
rect 23216 2148 23240 2150
rect 22920 2139 23296 2148
rect 28552 1170 28580 2314
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 28920 2204 29296 2213
rect 28976 2202 29000 2204
rect 29056 2202 29080 2204
rect 29136 2202 29160 2204
rect 29216 2202 29240 2204
rect 28976 2150 28986 2202
rect 29230 2150 29240 2202
rect 28976 2148 29000 2150
rect 29056 2148 29080 2150
rect 29136 2148 29160 2150
rect 29216 2148 29240 2150
rect 28920 2139 29296 2148
rect 30852 1465 30880 2246
rect 30838 1456 30894 1465
rect 30838 1391 30894 1400
rect 28368 1142 28580 1170
rect 28368 800 28396 1142
rect 18 0 74 800
rect 5170 0 5226 800
rect 10966 0 11022 800
rect 16762 0 16818 800
rect 22558 0 22614 800
rect 28354 0 28410 800
<< via2 >>
rect 4180 32122 4236 32124
rect 4260 32122 4316 32124
rect 4340 32122 4396 32124
rect 4420 32122 4476 32124
rect 4500 32122 4556 32124
rect 4180 32070 4182 32122
rect 4182 32070 4234 32122
rect 4234 32070 4236 32122
rect 4260 32070 4298 32122
rect 4298 32070 4310 32122
rect 4310 32070 4316 32122
rect 4340 32070 4362 32122
rect 4362 32070 4374 32122
rect 4374 32070 4396 32122
rect 4420 32070 4426 32122
rect 4426 32070 4438 32122
rect 4438 32070 4476 32122
rect 4500 32070 4502 32122
rect 4502 32070 4554 32122
rect 4554 32070 4556 32122
rect 4180 32068 4236 32070
rect 4260 32068 4316 32070
rect 4340 32068 4396 32070
rect 4420 32068 4476 32070
rect 4500 32068 4556 32070
rect 10180 32122 10236 32124
rect 10260 32122 10316 32124
rect 10340 32122 10396 32124
rect 10420 32122 10476 32124
rect 10500 32122 10556 32124
rect 10180 32070 10182 32122
rect 10182 32070 10234 32122
rect 10234 32070 10236 32122
rect 10260 32070 10298 32122
rect 10298 32070 10310 32122
rect 10310 32070 10316 32122
rect 10340 32070 10362 32122
rect 10362 32070 10374 32122
rect 10374 32070 10396 32122
rect 10420 32070 10426 32122
rect 10426 32070 10438 32122
rect 10438 32070 10476 32122
rect 10500 32070 10502 32122
rect 10502 32070 10554 32122
rect 10554 32070 10556 32122
rect 10180 32068 10236 32070
rect 10260 32068 10316 32070
rect 10340 32068 10396 32070
rect 10420 32068 10476 32070
rect 10500 32068 10556 32070
rect 16180 32122 16236 32124
rect 16260 32122 16316 32124
rect 16340 32122 16396 32124
rect 16420 32122 16476 32124
rect 16500 32122 16556 32124
rect 16180 32070 16182 32122
rect 16182 32070 16234 32122
rect 16234 32070 16236 32122
rect 16260 32070 16298 32122
rect 16298 32070 16310 32122
rect 16310 32070 16316 32122
rect 16340 32070 16362 32122
rect 16362 32070 16374 32122
rect 16374 32070 16396 32122
rect 16420 32070 16426 32122
rect 16426 32070 16438 32122
rect 16438 32070 16476 32122
rect 16500 32070 16502 32122
rect 16502 32070 16554 32122
rect 16554 32070 16556 32122
rect 16180 32068 16236 32070
rect 16260 32068 16316 32070
rect 16340 32068 16396 32070
rect 16420 32068 16476 32070
rect 16500 32068 16556 32070
rect 22180 32122 22236 32124
rect 22260 32122 22316 32124
rect 22340 32122 22396 32124
rect 22420 32122 22476 32124
rect 22500 32122 22556 32124
rect 22180 32070 22182 32122
rect 22182 32070 22234 32122
rect 22234 32070 22236 32122
rect 22260 32070 22298 32122
rect 22298 32070 22310 32122
rect 22310 32070 22316 32122
rect 22340 32070 22362 32122
rect 22362 32070 22374 32122
rect 22374 32070 22396 32122
rect 22420 32070 22426 32122
rect 22426 32070 22438 32122
rect 22438 32070 22476 32122
rect 22500 32070 22502 32122
rect 22502 32070 22554 32122
rect 22554 32070 22556 32122
rect 22180 32068 22236 32070
rect 22260 32068 22316 32070
rect 22340 32068 22396 32070
rect 22420 32068 22476 32070
rect 22500 32068 22556 32070
rect 28180 32122 28236 32124
rect 28260 32122 28316 32124
rect 28340 32122 28396 32124
rect 28420 32122 28476 32124
rect 28500 32122 28556 32124
rect 28180 32070 28182 32122
rect 28182 32070 28234 32122
rect 28234 32070 28236 32122
rect 28260 32070 28298 32122
rect 28298 32070 28310 32122
rect 28310 32070 28316 32122
rect 28340 32070 28362 32122
rect 28362 32070 28374 32122
rect 28374 32070 28396 32122
rect 28420 32070 28426 32122
rect 28426 32070 28438 32122
rect 28438 32070 28476 32122
rect 28500 32070 28502 32122
rect 28502 32070 28554 32122
rect 28554 32070 28556 32122
rect 28180 32068 28236 32070
rect 28260 32068 28316 32070
rect 28340 32068 28396 32070
rect 28420 32068 28476 32070
rect 28500 32068 28556 32070
rect 938 29960 994 30016
rect 938 23840 994 23896
rect 4920 31578 4976 31580
rect 5000 31578 5056 31580
rect 5080 31578 5136 31580
rect 5160 31578 5216 31580
rect 5240 31578 5296 31580
rect 4920 31526 4922 31578
rect 4922 31526 4974 31578
rect 4974 31526 4976 31578
rect 5000 31526 5038 31578
rect 5038 31526 5050 31578
rect 5050 31526 5056 31578
rect 5080 31526 5102 31578
rect 5102 31526 5114 31578
rect 5114 31526 5136 31578
rect 5160 31526 5166 31578
rect 5166 31526 5178 31578
rect 5178 31526 5216 31578
rect 5240 31526 5242 31578
rect 5242 31526 5294 31578
rect 5294 31526 5296 31578
rect 4920 31524 4976 31526
rect 5000 31524 5056 31526
rect 5080 31524 5136 31526
rect 5160 31524 5216 31526
rect 5240 31524 5296 31526
rect 10920 31578 10976 31580
rect 11000 31578 11056 31580
rect 11080 31578 11136 31580
rect 11160 31578 11216 31580
rect 11240 31578 11296 31580
rect 10920 31526 10922 31578
rect 10922 31526 10974 31578
rect 10974 31526 10976 31578
rect 11000 31526 11038 31578
rect 11038 31526 11050 31578
rect 11050 31526 11056 31578
rect 11080 31526 11102 31578
rect 11102 31526 11114 31578
rect 11114 31526 11136 31578
rect 11160 31526 11166 31578
rect 11166 31526 11178 31578
rect 11178 31526 11216 31578
rect 11240 31526 11242 31578
rect 11242 31526 11294 31578
rect 11294 31526 11296 31578
rect 10920 31524 10976 31526
rect 11000 31524 11056 31526
rect 11080 31524 11136 31526
rect 11160 31524 11216 31526
rect 11240 31524 11296 31526
rect 16920 31578 16976 31580
rect 17000 31578 17056 31580
rect 17080 31578 17136 31580
rect 17160 31578 17216 31580
rect 17240 31578 17296 31580
rect 16920 31526 16922 31578
rect 16922 31526 16974 31578
rect 16974 31526 16976 31578
rect 17000 31526 17038 31578
rect 17038 31526 17050 31578
rect 17050 31526 17056 31578
rect 17080 31526 17102 31578
rect 17102 31526 17114 31578
rect 17114 31526 17136 31578
rect 17160 31526 17166 31578
rect 17166 31526 17178 31578
rect 17178 31526 17216 31578
rect 17240 31526 17242 31578
rect 17242 31526 17294 31578
rect 17294 31526 17296 31578
rect 16920 31524 16976 31526
rect 17000 31524 17056 31526
rect 17080 31524 17136 31526
rect 17160 31524 17216 31526
rect 17240 31524 17296 31526
rect 4180 31034 4236 31036
rect 4260 31034 4316 31036
rect 4340 31034 4396 31036
rect 4420 31034 4476 31036
rect 4500 31034 4556 31036
rect 4180 30982 4182 31034
rect 4182 30982 4234 31034
rect 4234 30982 4236 31034
rect 4260 30982 4298 31034
rect 4298 30982 4310 31034
rect 4310 30982 4316 31034
rect 4340 30982 4362 31034
rect 4362 30982 4374 31034
rect 4374 30982 4396 31034
rect 4420 30982 4426 31034
rect 4426 30982 4438 31034
rect 4438 30982 4476 31034
rect 4500 30982 4502 31034
rect 4502 30982 4554 31034
rect 4554 30982 4556 31034
rect 4180 30980 4236 30982
rect 4260 30980 4316 30982
rect 4340 30980 4396 30982
rect 4420 30980 4476 30982
rect 4500 30980 4556 30982
rect 4920 30490 4976 30492
rect 5000 30490 5056 30492
rect 5080 30490 5136 30492
rect 5160 30490 5216 30492
rect 5240 30490 5296 30492
rect 4920 30438 4922 30490
rect 4922 30438 4974 30490
rect 4974 30438 4976 30490
rect 5000 30438 5038 30490
rect 5038 30438 5050 30490
rect 5050 30438 5056 30490
rect 5080 30438 5102 30490
rect 5102 30438 5114 30490
rect 5114 30438 5136 30490
rect 5160 30438 5166 30490
rect 5166 30438 5178 30490
rect 5178 30438 5216 30490
rect 5240 30438 5242 30490
rect 5242 30438 5294 30490
rect 5294 30438 5296 30490
rect 4920 30436 4976 30438
rect 5000 30436 5056 30438
rect 5080 30436 5136 30438
rect 5160 30436 5216 30438
rect 5240 30436 5296 30438
rect 4180 29946 4236 29948
rect 4260 29946 4316 29948
rect 4340 29946 4396 29948
rect 4420 29946 4476 29948
rect 4500 29946 4556 29948
rect 4180 29894 4182 29946
rect 4182 29894 4234 29946
rect 4234 29894 4236 29946
rect 4260 29894 4298 29946
rect 4298 29894 4310 29946
rect 4310 29894 4316 29946
rect 4340 29894 4362 29946
rect 4362 29894 4374 29946
rect 4374 29894 4396 29946
rect 4420 29894 4426 29946
rect 4426 29894 4438 29946
rect 4438 29894 4476 29946
rect 4500 29894 4502 29946
rect 4502 29894 4554 29946
rect 4554 29894 4556 29946
rect 4180 29892 4236 29894
rect 4260 29892 4316 29894
rect 4340 29892 4396 29894
rect 4420 29892 4476 29894
rect 4500 29892 4556 29894
rect 4920 29402 4976 29404
rect 5000 29402 5056 29404
rect 5080 29402 5136 29404
rect 5160 29402 5216 29404
rect 5240 29402 5296 29404
rect 4920 29350 4922 29402
rect 4922 29350 4974 29402
rect 4974 29350 4976 29402
rect 5000 29350 5038 29402
rect 5038 29350 5050 29402
rect 5050 29350 5056 29402
rect 5080 29350 5102 29402
rect 5102 29350 5114 29402
rect 5114 29350 5136 29402
rect 5160 29350 5166 29402
rect 5166 29350 5178 29402
rect 5178 29350 5216 29402
rect 5240 29350 5242 29402
rect 5242 29350 5294 29402
rect 5294 29350 5296 29402
rect 4920 29348 4976 29350
rect 5000 29348 5056 29350
rect 5080 29348 5136 29350
rect 5160 29348 5216 29350
rect 5240 29348 5296 29350
rect 4180 28858 4236 28860
rect 4260 28858 4316 28860
rect 4340 28858 4396 28860
rect 4420 28858 4476 28860
rect 4500 28858 4556 28860
rect 4180 28806 4182 28858
rect 4182 28806 4234 28858
rect 4234 28806 4236 28858
rect 4260 28806 4298 28858
rect 4298 28806 4310 28858
rect 4310 28806 4316 28858
rect 4340 28806 4362 28858
rect 4362 28806 4374 28858
rect 4374 28806 4396 28858
rect 4420 28806 4426 28858
rect 4426 28806 4438 28858
rect 4438 28806 4476 28858
rect 4500 28806 4502 28858
rect 4502 28806 4554 28858
rect 4554 28806 4556 28858
rect 4180 28804 4236 28806
rect 4260 28804 4316 28806
rect 4340 28804 4396 28806
rect 4420 28804 4476 28806
rect 4500 28804 4556 28806
rect 4920 28314 4976 28316
rect 5000 28314 5056 28316
rect 5080 28314 5136 28316
rect 5160 28314 5216 28316
rect 5240 28314 5296 28316
rect 4920 28262 4922 28314
rect 4922 28262 4974 28314
rect 4974 28262 4976 28314
rect 5000 28262 5038 28314
rect 5038 28262 5050 28314
rect 5050 28262 5056 28314
rect 5080 28262 5102 28314
rect 5102 28262 5114 28314
rect 5114 28262 5136 28314
rect 5160 28262 5166 28314
rect 5166 28262 5178 28314
rect 5178 28262 5216 28314
rect 5240 28262 5242 28314
rect 5242 28262 5294 28314
rect 5294 28262 5296 28314
rect 4920 28260 4976 28262
rect 5000 28260 5056 28262
rect 5080 28260 5136 28262
rect 5160 28260 5216 28262
rect 5240 28260 5296 28262
rect 4180 27770 4236 27772
rect 4260 27770 4316 27772
rect 4340 27770 4396 27772
rect 4420 27770 4476 27772
rect 4500 27770 4556 27772
rect 4180 27718 4182 27770
rect 4182 27718 4234 27770
rect 4234 27718 4236 27770
rect 4260 27718 4298 27770
rect 4298 27718 4310 27770
rect 4310 27718 4316 27770
rect 4340 27718 4362 27770
rect 4362 27718 4374 27770
rect 4374 27718 4396 27770
rect 4420 27718 4426 27770
rect 4426 27718 4438 27770
rect 4438 27718 4476 27770
rect 4500 27718 4502 27770
rect 4502 27718 4554 27770
rect 4554 27718 4556 27770
rect 4180 27716 4236 27718
rect 4260 27716 4316 27718
rect 4340 27716 4396 27718
rect 4420 27716 4476 27718
rect 4500 27716 4556 27718
rect 10180 31034 10236 31036
rect 10260 31034 10316 31036
rect 10340 31034 10396 31036
rect 10420 31034 10476 31036
rect 10500 31034 10556 31036
rect 10180 30982 10182 31034
rect 10182 30982 10234 31034
rect 10234 30982 10236 31034
rect 10260 30982 10298 31034
rect 10298 30982 10310 31034
rect 10310 30982 10316 31034
rect 10340 30982 10362 31034
rect 10362 30982 10374 31034
rect 10374 30982 10396 31034
rect 10420 30982 10426 31034
rect 10426 30982 10438 31034
rect 10438 30982 10476 31034
rect 10500 30982 10502 31034
rect 10502 30982 10554 31034
rect 10554 30982 10556 31034
rect 10180 30980 10236 30982
rect 10260 30980 10316 30982
rect 10340 30980 10396 30982
rect 10420 30980 10476 30982
rect 10500 30980 10556 30982
rect 4920 27226 4976 27228
rect 5000 27226 5056 27228
rect 5080 27226 5136 27228
rect 5160 27226 5216 27228
rect 5240 27226 5296 27228
rect 4920 27174 4922 27226
rect 4922 27174 4974 27226
rect 4974 27174 4976 27226
rect 5000 27174 5038 27226
rect 5038 27174 5050 27226
rect 5050 27174 5056 27226
rect 5080 27174 5102 27226
rect 5102 27174 5114 27226
rect 5114 27174 5136 27226
rect 5160 27174 5166 27226
rect 5166 27174 5178 27226
rect 5178 27174 5216 27226
rect 5240 27174 5242 27226
rect 5242 27174 5294 27226
rect 5294 27174 5296 27226
rect 4920 27172 4976 27174
rect 5000 27172 5056 27174
rect 5080 27172 5136 27174
rect 5160 27172 5216 27174
rect 5240 27172 5296 27174
rect 4180 26682 4236 26684
rect 4260 26682 4316 26684
rect 4340 26682 4396 26684
rect 4420 26682 4476 26684
rect 4500 26682 4556 26684
rect 4180 26630 4182 26682
rect 4182 26630 4234 26682
rect 4234 26630 4236 26682
rect 4260 26630 4298 26682
rect 4298 26630 4310 26682
rect 4310 26630 4316 26682
rect 4340 26630 4362 26682
rect 4362 26630 4374 26682
rect 4374 26630 4396 26682
rect 4420 26630 4426 26682
rect 4426 26630 4438 26682
rect 4438 26630 4476 26682
rect 4500 26630 4502 26682
rect 4502 26630 4554 26682
rect 4554 26630 4556 26682
rect 4180 26628 4236 26630
rect 4260 26628 4316 26630
rect 4340 26628 4396 26630
rect 4420 26628 4476 26630
rect 4500 26628 4556 26630
rect 4920 26138 4976 26140
rect 5000 26138 5056 26140
rect 5080 26138 5136 26140
rect 5160 26138 5216 26140
rect 5240 26138 5296 26140
rect 4920 26086 4922 26138
rect 4922 26086 4974 26138
rect 4974 26086 4976 26138
rect 5000 26086 5038 26138
rect 5038 26086 5050 26138
rect 5050 26086 5056 26138
rect 5080 26086 5102 26138
rect 5102 26086 5114 26138
rect 5114 26086 5136 26138
rect 5160 26086 5166 26138
rect 5166 26086 5178 26138
rect 5178 26086 5216 26138
rect 5240 26086 5242 26138
rect 5242 26086 5294 26138
rect 5294 26086 5296 26138
rect 4920 26084 4976 26086
rect 5000 26084 5056 26086
rect 5080 26084 5136 26086
rect 5160 26084 5216 26086
rect 5240 26084 5296 26086
rect 4180 25594 4236 25596
rect 4260 25594 4316 25596
rect 4340 25594 4396 25596
rect 4420 25594 4476 25596
rect 4500 25594 4556 25596
rect 4180 25542 4182 25594
rect 4182 25542 4234 25594
rect 4234 25542 4236 25594
rect 4260 25542 4298 25594
rect 4298 25542 4310 25594
rect 4310 25542 4316 25594
rect 4340 25542 4362 25594
rect 4362 25542 4374 25594
rect 4374 25542 4396 25594
rect 4420 25542 4426 25594
rect 4426 25542 4438 25594
rect 4438 25542 4476 25594
rect 4500 25542 4502 25594
rect 4502 25542 4554 25594
rect 4554 25542 4556 25594
rect 4180 25540 4236 25542
rect 4260 25540 4316 25542
rect 4340 25540 4396 25542
rect 4420 25540 4476 25542
rect 4500 25540 4556 25542
rect 4180 24506 4236 24508
rect 4260 24506 4316 24508
rect 4340 24506 4396 24508
rect 4420 24506 4476 24508
rect 4500 24506 4556 24508
rect 4180 24454 4182 24506
rect 4182 24454 4234 24506
rect 4234 24454 4236 24506
rect 4260 24454 4298 24506
rect 4298 24454 4310 24506
rect 4310 24454 4316 24506
rect 4340 24454 4362 24506
rect 4362 24454 4374 24506
rect 4374 24454 4396 24506
rect 4420 24454 4426 24506
rect 4426 24454 4438 24506
rect 4438 24454 4476 24506
rect 4500 24454 4502 24506
rect 4502 24454 4554 24506
rect 4554 24454 4556 24506
rect 4180 24452 4236 24454
rect 4260 24452 4316 24454
rect 4340 24452 4396 24454
rect 4420 24452 4476 24454
rect 4500 24452 4556 24454
rect 4180 23418 4236 23420
rect 4260 23418 4316 23420
rect 4340 23418 4396 23420
rect 4420 23418 4476 23420
rect 4500 23418 4556 23420
rect 4180 23366 4182 23418
rect 4182 23366 4234 23418
rect 4234 23366 4236 23418
rect 4260 23366 4298 23418
rect 4298 23366 4310 23418
rect 4310 23366 4316 23418
rect 4340 23366 4362 23418
rect 4362 23366 4374 23418
rect 4374 23366 4396 23418
rect 4420 23366 4426 23418
rect 4426 23366 4438 23418
rect 4438 23366 4476 23418
rect 4500 23366 4502 23418
rect 4502 23366 4554 23418
rect 4554 23366 4556 23418
rect 4180 23364 4236 23366
rect 4260 23364 4316 23366
rect 4340 23364 4396 23366
rect 4420 23364 4476 23366
rect 4500 23364 4556 23366
rect 4920 25050 4976 25052
rect 5000 25050 5056 25052
rect 5080 25050 5136 25052
rect 5160 25050 5216 25052
rect 5240 25050 5296 25052
rect 4920 24998 4922 25050
rect 4922 24998 4974 25050
rect 4974 24998 4976 25050
rect 5000 24998 5038 25050
rect 5038 24998 5050 25050
rect 5050 24998 5056 25050
rect 5080 24998 5102 25050
rect 5102 24998 5114 25050
rect 5114 24998 5136 25050
rect 5160 24998 5166 25050
rect 5166 24998 5178 25050
rect 5178 24998 5216 25050
rect 5240 24998 5242 25050
rect 5242 24998 5294 25050
rect 5294 24998 5296 25050
rect 4920 24996 4976 24998
rect 5000 24996 5056 24998
rect 5080 24996 5136 24998
rect 5160 24996 5216 24998
rect 5240 24996 5296 24998
rect 4180 22330 4236 22332
rect 4260 22330 4316 22332
rect 4340 22330 4396 22332
rect 4420 22330 4476 22332
rect 4500 22330 4556 22332
rect 4180 22278 4182 22330
rect 4182 22278 4234 22330
rect 4234 22278 4236 22330
rect 4260 22278 4298 22330
rect 4298 22278 4310 22330
rect 4310 22278 4316 22330
rect 4340 22278 4362 22330
rect 4362 22278 4374 22330
rect 4374 22278 4396 22330
rect 4420 22278 4426 22330
rect 4426 22278 4438 22330
rect 4438 22278 4476 22330
rect 4500 22278 4502 22330
rect 4502 22278 4554 22330
rect 4554 22278 4556 22330
rect 4180 22276 4236 22278
rect 4260 22276 4316 22278
rect 4340 22276 4396 22278
rect 4420 22276 4476 22278
rect 4500 22276 4556 22278
rect 4920 23962 4976 23964
rect 5000 23962 5056 23964
rect 5080 23962 5136 23964
rect 5160 23962 5216 23964
rect 5240 23962 5296 23964
rect 4920 23910 4922 23962
rect 4922 23910 4974 23962
rect 4974 23910 4976 23962
rect 5000 23910 5038 23962
rect 5038 23910 5050 23962
rect 5050 23910 5056 23962
rect 5080 23910 5102 23962
rect 5102 23910 5114 23962
rect 5114 23910 5136 23962
rect 5160 23910 5166 23962
rect 5166 23910 5178 23962
rect 5178 23910 5216 23962
rect 5240 23910 5242 23962
rect 5242 23910 5294 23962
rect 5294 23910 5296 23962
rect 4920 23908 4976 23910
rect 5000 23908 5056 23910
rect 5080 23908 5136 23910
rect 5160 23908 5216 23910
rect 5240 23908 5296 23910
rect 4920 22874 4976 22876
rect 5000 22874 5056 22876
rect 5080 22874 5136 22876
rect 5160 22874 5216 22876
rect 5240 22874 5296 22876
rect 4920 22822 4922 22874
rect 4922 22822 4974 22874
rect 4974 22822 4976 22874
rect 5000 22822 5038 22874
rect 5038 22822 5050 22874
rect 5050 22822 5056 22874
rect 5080 22822 5102 22874
rect 5102 22822 5114 22874
rect 5114 22822 5136 22874
rect 5160 22822 5166 22874
rect 5166 22822 5178 22874
rect 5178 22822 5216 22874
rect 5240 22822 5242 22874
rect 5242 22822 5294 22874
rect 5294 22822 5296 22874
rect 4920 22820 4976 22822
rect 5000 22820 5056 22822
rect 5080 22820 5136 22822
rect 5160 22820 5216 22822
rect 5240 22820 5296 22822
rect 4180 21242 4236 21244
rect 4260 21242 4316 21244
rect 4340 21242 4396 21244
rect 4420 21242 4476 21244
rect 4500 21242 4556 21244
rect 4180 21190 4182 21242
rect 4182 21190 4234 21242
rect 4234 21190 4236 21242
rect 4260 21190 4298 21242
rect 4298 21190 4310 21242
rect 4310 21190 4316 21242
rect 4340 21190 4362 21242
rect 4362 21190 4374 21242
rect 4374 21190 4396 21242
rect 4420 21190 4426 21242
rect 4426 21190 4438 21242
rect 4438 21190 4476 21242
rect 4500 21190 4502 21242
rect 4502 21190 4554 21242
rect 4554 21190 4556 21242
rect 4180 21188 4236 21190
rect 4260 21188 4316 21190
rect 4340 21188 4396 21190
rect 4420 21188 4476 21190
rect 4500 21188 4556 21190
rect 4180 20154 4236 20156
rect 4260 20154 4316 20156
rect 4340 20154 4396 20156
rect 4420 20154 4476 20156
rect 4500 20154 4556 20156
rect 4180 20102 4182 20154
rect 4182 20102 4234 20154
rect 4234 20102 4236 20154
rect 4260 20102 4298 20154
rect 4298 20102 4310 20154
rect 4310 20102 4316 20154
rect 4340 20102 4362 20154
rect 4362 20102 4374 20154
rect 4374 20102 4396 20154
rect 4420 20102 4426 20154
rect 4426 20102 4438 20154
rect 4438 20102 4476 20154
rect 4500 20102 4502 20154
rect 4502 20102 4554 20154
rect 4554 20102 4556 20154
rect 4180 20100 4236 20102
rect 4260 20100 4316 20102
rect 4340 20100 4396 20102
rect 4420 20100 4476 20102
rect 4500 20100 4556 20102
rect 1398 17856 1454 17912
rect 4180 19066 4236 19068
rect 4260 19066 4316 19068
rect 4340 19066 4396 19068
rect 4420 19066 4476 19068
rect 4500 19066 4556 19068
rect 4180 19014 4182 19066
rect 4182 19014 4234 19066
rect 4234 19014 4236 19066
rect 4260 19014 4298 19066
rect 4298 19014 4310 19066
rect 4310 19014 4316 19066
rect 4340 19014 4362 19066
rect 4362 19014 4374 19066
rect 4374 19014 4396 19066
rect 4420 19014 4426 19066
rect 4426 19014 4438 19066
rect 4438 19014 4476 19066
rect 4500 19014 4502 19066
rect 4502 19014 4554 19066
rect 4554 19014 4556 19066
rect 4180 19012 4236 19014
rect 4260 19012 4316 19014
rect 4340 19012 4396 19014
rect 4420 19012 4476 19014
rect 4500 19012 4556 19014
rect 4920 21786 4976 21788
rect 5000 21786 5056 21788
rect 5080 21786 5136 21788
rect 5160 21786 5216 21788
rect 5240 21786 5296 21788
rect 4920 21734 4922 21786
rect 4922 21734 4974 21786
rect 4974 21734 4976 21786
rect 5000 21734 5038 21786
rect 5038 21734 5050 21786
rect 5050 21734 5056 21786
rect 5080 21734 5102 21786
rect 5102 21734 5114 21786
rect 5114 21734 5136 21786
rect 5160 21734 5166 21786
rect 5166 21734 5178 21786
rect 5178 21734 5216 21786
rect 5240 21734 5242 21786
rect 5242 21734 5294 21786
rect 5294 21734 5296 21786
rect 4920 21732 4976 21734
rect 5000 21732 5056 21734
rect 5080 21732 5136 21734
rect 5160 21732 5216 21734
rect 5240 21732 5296 21734
rect 4920 20698 4976 20700
rect 5000 20698 5056 20700
rect 5080 20698 5136 20700
rect 5160 20698 5216 20700
rect 5240 20698 5296 20700
rect 4920 20646 4922 20698
rect 4922 20646 4974 20698
rect 4974 20646 4976 20698
rect 5000 20646 5038 20698
rect 5038 20646 5050 20698
rect 5050 20646 5056 20698
rect 5080 20646 5102 20698
rect 5102 20646 5114 20698
rect 5114 20646 5136 20698
rect 5160 20646 5166 20698
rect 5166 20646 5178 20698
rect 5178 20646 5216 20698
rect 5240 20646 5242 20698
rect 5242 20646 5294 20698
rect 5294 20646 5296 20698
rect 4920 20644 4976 20646
rect 5000 20644 5056 20646
rect 5080 20644 5136 20646
rect 5160 20644 5216 20646
rect 5240 20644 5296 20646
rect 4920 19610 4976 19612
rect 5000 19610 5056 19612
rect 5080 19610 5136 19612
rect 5160 19610 5216 19612
rect 5240 19610 5296 19612
rect 4920 19558 4922 19610
rect 4922 19558 4974 19610
rect 4974 19558 4976 19610
rect 5000 19558 5038 19610
rect 5038 19558 5050 19610
rect 5050 19558 5056 19610
rect 5080 19558 5102 19610
rect 5102 19558 5114 19610
rect 5114 19558 5136 19610
rect 5160 19558 5166 19610
rect 5166 19558 5178 19610
rect 5178 19558 5216 19610
rect 5240 19558 5242 19610
rect 5242 19558 5294 19610
rect 5294 19558 5296 19610
rect 4920 19556 4976 19558
rect 5000 19556 5056 19558
rect 5080 19556 5136 19558
rect 5160 19556 5216 19558
rect 5240 19556 5296 19558
rect 4180 17978 4236 17980
rect 4260 17978 4316 17980
rect 4340 17978 4396 17980
rect 4420 17978 4476 17980
rect 4500 17978 4556 17980
rect 4180 17926 4182 17978
rect 4182 17926 4234 17978
rect 4234 17926 4236 17978
rect 4260 17926 4298 17978
rect 4298 17926 4310 17978
rect 4310 17926 4316 17978
rect 4340 17926 4362 17978
rect 4362 17926 4374 17978
rect 4374 17926 4396 17978
rect 4420 17926 4426 17978
rect 4426 17926 4438 17978
rect 4438 17926 4476 17978
rect 4500 17926 4502 17978
rect 4502 17926 4554 17978
rect 4554 17926 4556 17978
rect 4180 17924 4236 17926
rect 4260 17924 4316 17926
rect 4340 17924 4396 17926
rect 4420 17924 4476 17926
rect 4500 17924 4556 17926
rect 4180 16890 4236 16892
rect 4260 16890 4316 16892
rect 4340 16890 4396 16892
rect 4420 16890 4476 16892
rect 4500 16890 4556 16892
rect 4180 16838 4182 16890
rect 4182 16838 4234 16890
rect 4234 16838 4236 16890
rect 4260 16838 4298 16890
rect 4298 16838 4310 16890
rect 4310 16838 4316 16890
rect 4340 16838 4362 16890
rect 4362 16838 4374 16890
rect 4374 16838 4396 16890
rect 4420 16838 4426 16890
rect 4426 16838 4438 16890
rect 4438 16838 4476 16890
rect 4500 16838 4502 16890
rect 4502 16838 4554 16890
rect 4554 16838 4556 16890
rect 4180 16836 4236 16838
rect 4260 16836 4316 16838
rect 4340 16836 4396 16838
rect 4420 16836 4476 16838
rect 4500 16836 4556 16838
rect 4180 15802 4236 15804
rect 4260 15802 4316 15804
rect 4340 15802 4396 15804
rect 4420 15802 4476 15804
rect 4500 15802 4556 15804
rect 4180 15750 4182 15802
rect 4182 15750 4234 15802
rect 4234 15750 4236 15802
rect 4260 15750 4298 15802
rect 4298 15750 4310 15802
rect 4310 15750 4316 15802
rect 4340 15750 4362 15802
rect 4362 15750 4374 15802
rect 4374 15750 4396 15802
rect 4420 15750 4426 15802
rect 4426 15750 4438 15802
rect 4438 15750 4476 15802
rect 4500 15750 4502 15802
rect 4502 15750 4554 15802
rect 4554 15750 4556 15802
rect 4180 15748 4236 15750
rect 4260 15748 4316 15750
rect 4340 15748 4396 15750
rect 4420 15748 4476 15750
rect 4500 15748 4556 15750
rect 4180 14714 4236 14716
rect 4260 14714 4316 14716
rect 4340 14714 4396 14716
rect 4420 14714 4476 14716
rect 4500 14714 4556 14716
rect 4180 14662 4182 14714
rect 4182 14662 4234 14714
rect 4234 14662 4236 14714
rect 4260 14662 4298 14714
rect 4298 14662 4310 14714
rect 4310 14662 4316 14714
rect 4340 14662 4362 14714
rect 4362 14662 4374 14714
rect 4374 14662 4396 14714
rect 4420 14662 4426 14714
rect 4426 14662 4438 14714
rect 4438 14662 4476 14714
rect 4500 14662 4502 14714
rect 4502 14662 4554 14714
rect 4554 14662 4556 14714
rect 4180 14660 4236 14662
rect 4260 14660 4316 14662
rect 4340 14660 4396 14662
rect 4420 14660 4476 14662
rect 4500 14660 4556 14662
rect 938 11600 994 11656
rect 4180 13626 4236 13628
rect 4260 13626 4316 13628
rect 4340 13626 4396 13628
rect 4420 13626 4476 13628
rect 4500 13626 4556 13628
rect 4180 13574 4182 13626
rect 4182 13574 4234 13626
rect 4234 13574 4236 13626
rect 4260 13574 4298 13626
rect 4298 13574 4310 13626
rect 4310 13574 4316 13626
rect 4340 13574 4362 13626
rect 4362 13574 4374 13626
rect 4374 13574 4396 13626
rect 4420 13574 4426 13626
rect 4426 13574 4438 13626
rect 4438 13574 4476 13626
rect 4500 13574 4502 13626
rect 4502 13574 4554 13626
rect 4554 13574 4556 13626
rect 4180 13572 4236 13574
rect 4260 13572 4316 13574
rect 4340 13572 4396 13574
rect 4420 13572 4476 13574
rect 4500 13572 4556 13574
rect 4920 18522 4976 18524
rect 5000 18522 5056 18524
rect 5080 18522 5136 18524
rect 5160 18522 5216 18524
rect 5240 18522 5296 18524
rect 4920 18470 4922 18522
rect 4922 18470 4974 18522
rect 4974 18470 4976 18522
rect 5000 18470 5038 18522
rect 5038 18470 5050 18522
rect 5050 18470 5056 18522
rect 5080 18470 5102 18522
rect 5102 18470 5114 18522
rect 5114 18470 5136 18522
rect 5160 18470 5166 18522
rect 5166 18470 5178 18522
rect 5178 18470 5216 18522
rect 5240 18470 5242 18522
rect 5242 18470 5294 18522
rect 5294 18470 5296 18522
rect 4920 18468 4976 18470
rect 5000 18468 5056 18470
rect 5080 18468 5136 18470
rect 5160 18468 5216 18470
rect 5240 18468 5296 18470
rect 4920 17434 4976 17436
rect 5000 17434 5056 17436
rect 5080 17434 5136 17436
rect 5160 17434 5216 17436
rect 5240 17434 5296 17436
rect 4920 17382 4922 17434
rect 4922 17382 4974 17434
rect 4974 17382 4976 17434
rect 5000 17382 5038 17434
rect 5038 17382 5050 17434
rect 5050 17382 5056 17434
rect 5080 17382 5102 17434
rect 5102 17382 5114 17434
rect 5114 17382 5136 17434
rect 5160 17382 5166 17434
rect 5166 17382 5178 17434
rect 5178 17382 5216 17434
rect 5240 17382 5242 17434
rect 5242 17382 5294 17434
rect 5294 17382 5296 17434
rect 4920 17380 4976 17382
rect 5000 17380 5056 17382
rect 5080 17380 5136 17382
rect 5160 17380 5216 17382
rect 5240 17380 5296 17382
rect 4920 16346 4976 16348
rect 5000 16346 5056 16348
rect 5080 16346 5136 16348
rect 5160 16346 5216 16348
rect 5240 16346 5296 16348
rect 4920 16294 4922 16346
rect 4922 16294 4974 16346
rect 4974 16294 4976 16346
rect 5000 16294 5038 16346
rect 5038 16294 5050 16346
rect 5050 16294 5056 16346
rect 5080 16294 5102 16346
rect 5102 16294 5114 16346
rect 5114 16294 5136 16346
rect 5160 16294 5166 16346
rect 5166 16294 5178 16346
rect 5178 16294 5216 16346
rect 5240 16294 5242 16346
rect 5242 16294 5294 16346
rect 5294 16294 5296 16346
rect 4920 16292 4976 16294
rect 5000 16292 5056 16294
rect 5080 16292 5136 16294
rect 5160 16292 5216 16294
rect 5240 16292 5296 16294
rect 4920 15258 4976 15260
rect 5000 15258 5056 15260
rect 5080 15258 5136 15260
rect 5160 15258 5216 15260
rect 5240 15258 5296 15260
rect 4920 15206 4922 15258
rect 4922 15206 4974 15258
rect 4974 15206 4976 15258
rect 5000 15206 5038 15258
rect 5038 15206 5050 15258
rect 5050 15206 5056 15258
rect 5080 15206 5102 15258
rect 5102 15206 5114 15258
rect 5114 15206 5136 15258
rect 5160 15206 5166 15258
rect 5166 15206 5178 15258
rect 5178 15206 5216 15258
rect 5240 15206 5242 15258
rect 5242 15206 5294 15258
rect 5294 15206 5296 15258
rect 4920 15204 4976 15206
rect 5000 15204 5056 15206
rect 5080 15204 5136 15206
rect 5160 15204 5216 15206
rect 5240 15204 5296 15206
rect 4920 14170 4976 14172
rect 5000 14170 5056 14172
rect 5080 14170 5136 14172
rect 5160 14170 5216 14172
rect 5240 14170 5296 14172
rect 4920 14118 4922 14170
rect 4922 14118 4974 14170
rect 4974 14118 4976 14170
rect 5000 14118 5038 14170
rect 5038 14118 5050 14170
rect 5050 14118 5056 14170
rect 5080 14118 5102 14170
rect 5102 14118 5114 14170
rect 5114 14118 5136 14170
rect 5160 14118 5166 14170
rect 5166 14118 5178 14170
rect 5178 14118 5216 14170
rect 5240 14118 5242 14170
rect 5242 14118 5294 14170
rect 5294 14118 5296 14170
rect 4920 14116 4976 14118
rect 5000 14116 5056 14118
rect 5080 14116 5136 14118
rect 5160 14116 5216 14118
rect 5240 14116 5296 14118
rect 4920 13082 4976 13084
rect 5000 13082 5056 13084
rect 5080 13082 5136 13084
rect 5160 13082 5216 13084
rect 5240 13082 5296 13084
rect 4920 13030 4922 13082
rect 4922 13030 4974 13082
rect 4974 13030 4976 13082
rect 5000 13030 5038 13082
rect 5038 13030 5050 13082
rect 5050 13030 5056 13082
rect 5080 13030 5102 13082
rect 5102 13030 5114 13082
rect 5114 13030 5136 13082
rect 5160 13030 5166 13082
rect 5166 13030 5178 13082
rect 5178 13030 5216 13082
rect 5240 13030 5242 13082
rect 5242 13030 5294 13082
rect 5294 13030 5296 13082
rect 4920 13028 4976 13030
rect 5000 13028 5056 13030
rect 5080 13028 5136 13030
rect 5160 13028 5216 13030
rect 5240 13028 5296 13030
rect 4180 12538 4236 12540
rect 4260 12538 4316 12540
rect 4340 12538 4396 12540
rect 4420 12538 4476 12540
rect 4500 12538 4556 12540
rect 4180 12486 4182 12538
rect 4182 12486 4234 12538
rect 4234 12486 4236 12538
rect 4260 12486 4298 12538
rect 4298 12486 4310 12538
rect 4310 12486 4316 12538
rect 4340 12486 4362 12538
rect 4362 12486 4374 12538
rect 4374 12486 4396 12538
rect 4420 12486 4426 12538
rect 4426 12486 4438 12538
rect 4438 12486 4476 12538
rect 4500 12486 4502 12538
rect 4502 12486 4554 12538
rect 4554 12486 4556 12538
rect 4180 12484 4236 12486
rect 4260 12484 4316 12486
rect 4340 12484 4396 12486
rect 4420 12484 4476 12486
rect 4500 12484 4556 12486
rect 4180 11450 4236 11452
rect 4260 11450 4316 11452
rect 4340 11450 4396 11452
rect 4420 11450 4476 11452
rect 4500 11450 4556 11452
rect 4180 11398 4182 11450
rect 4182 11398 4234 11450
rect 4234 11398 4236 11450
rect 4260 11398 4298 11450
rect 4298 11398 4310 11450
rect 4310 11398 4316 11450
rect 4340 11398 4362 11450
rect 4362 11398 4374 11450
rect 4374 11398 4396 11450
rect 4420 11398 4426 11450
rect 4426 11398 4438 11450
rect 4438 11398 4476 11450
rect 4500 11398 4502 11450
rect 4502 11398 4554 11450
rect 4554 11398 4556 11450
rect 4180 11396 4236 11398
rect 4260 11396 4316 11398
rect 4340 11396 4396 11398
rect 4420 11396 4476 11398
rect 4500 11396 4556 11398
rect 4920 11994 4976 11996
rect 5000 11994 5056 11996
rect 5080 11994 5136 11996
rect 5160 11994 5216 11996
rect 5240 11994 5296 11996
rect 4920 11942 4922 11994
rect 4922 11942 4974 11994
rect 4974 11942 4976 11994
rect 5000 11942 5038 11994
rect 5038 11942 5050 11994
rect 5050 11942 5056 11994
rect 5080 11942 5102 11994
rect 5102 11942 5114 11994
rect 5114 11942 5136 11994
rect 5160 11942 5166 11994
rect 5166 11942 5178 11994
rect 5178 11942 5216 11994
rect 5240 11942 5242 11994
rect 5242 11942 5294 11994
rect 5294 11942 5296 11994
rect 4920 11940 4976 11942
rect 5000 11940 5056 11942
rect 5080 11940 5136 11942
rect 5160 11940 5216 11942
rect 5240 11940 5296 11942
rect 4180 10362 4236 10364
rect 4260 10362 4316 10364
rect 4340 10362 4396 10364
rect 4420 10362 4476 10364
rect 4500 10362 4556 10364
rect 4180 10310 4182 10362
rect 4182 10310 4234 10362
rect 4234 10310 4236 10362
rect 4260 10310 4298 10362
rect 4298 10310 4310 10362
rect 4310 10310 4316 10362
rect 4340 10310 4362 10362
rect 4362 10310 4374 10362
rect 4374 10310 4396 10362
rect 4420 10310 4426 10362
rect 4426 10310 4438 10362
rect 4438 10310 4476 10362
rect 4500 10310 4502 10362
rect 4502 10310 4554 10362
rect 4554 10310 4556 10362
rect 4180 10308 4236 10310
rect 4260 10308 4316 10310
rect 4340 10308 4396 10310
rect 4420 10308 4476 10310
rect 4500 10308 4556 10310
rect 4920 10906 4976 10908
rect 5000 10906 5056 10908
rect 5080 10906 5136 10908
rect 5160 10906 5216 10908
rect 5240 10906 5296 10908
rect 4920 10854 4922 10906
rect 4922 10854 4974 10906
rect 4974 10854 4976 10906
rect 5000 10854 5038 10906
rect 5038 10854 5050 10906
rect 5050 10854 5056 10906
rect 5080 10854 5102 10906
rect 5102 10854 5114 10906
rect 5114 10854 5136 10906
rect 5160 10854 5166 10906
rect 5166 10854 5178 10906
rect 5178 10854 5216 10906
rect 5240 10854 5242 10906
rect 5242 10854 5294 10906
rect 5294 10854 5296 10906
rect 4920 10852 4976 10854
rect 5000 10852 5056 10854
rect 5080 10852 5136 10854
rect 5160 10852 5216 10854
rect 5240 10852 5296 10854
rect 4180 9274 4236 9276
rect 4260 9274 4316 9276
rect 4340 9274 4396 9276
rect 4420 9274 4476 9276
rect 4500 9274 4556 9276
rect 4180 9222 4182 9274
rect 4182 9222 4234 9274
rect 4234 9222 4236 9274
rect 4260 9222 4298 9274
rect 4298 9222 4310 9274
rect 4310 9222 4316 9274
rect 4340 9222 4362 9274
rect 4362 9222 4374 9274
rect 4374 9222 4396 9274
rect 4420 9222 4426 9274
rect 4426 9222 4438 9274
rect 4438 9222 4476 9274
rect 4500 9222 4502 9274
rect 4502 9222 4554 9274
rect 4554 9222 4556 9274
rect 4180 9220 4236 9222
rect 4260 9220 4316 9222
rect 4340 9220 4396 9222
rect 4420 9220 4476 9222
rect 4500 9220 4556 9222
rect 4920 9818 4976 9820
rect 5000 9818 5056 9820
rect 5080 9818 5136 9820
rect 5160 9818 5216 9820
rect 5240 9818 5296 9820
rect 4920 9766 4922 9818
rect 4922 9766 4974 9818
rect 4974 9766 4976 9818
rect 5000 9766 5038 9818
rect 5038 9766 5050 9818
rect 5050 9766 5056 9818
rect 5080 9766 5102 9818
rect 5102 9766 5114 9818
rect 5114 9766 5136 9818
rect 5160 9766 5166 9818
rect 5166 9766 5178 9818
rect 5178 9766 5216 9818
rect 5240 9766 5242 9818
rect 5242 9766 5294 9818
rect 5294 9766 5296 9818
rect 4920 9764 4976 9766
rect 5000 9764 5056 9766
rect 5080 9764 5136 9766
rect 5160 9764 5216 9766
rect 5240 9764 5296 9766
rect 4920 8730 4976 8732
rect 5000 8730 5056 8732
rect 5080 8730 5136 8732
rect 5160 8730 5216 8732
rect 5240 8730 5296 8732
rect 4920 8678 4922 8730
rect 4922 8678 4974 8730
rect 4974 8678 4976 8730
rect 5000 8678 5038 8730
rect 5038 8678 5050 8730
rect 5050 8678 5056 8730
rect 5080 8678 5102 8730
rect 5102 8678 5114 8730
rect 5114 8678 5136 8730
rect 5160 8678 5166 8730
rect 5166 8678 5178 8730
rect 5178 8678 5216 8730
rect 5240 8678 5242 8730
rect 5242 8678 5294 8730
rect 5294 8678 5296 8730
rect 4920 8676 4976 8678
rect 5000 8676 5056 8678
rect 5080 8676 5136 8678
rect 5160 8676 5216 8678
rect 5240 8676 5296 8678
rect 10920 30490 10976 30492
rect 11000 30490 11056 30492
rect 11080 30490 11136 30492
rect 11160 30490 11216 30492
rect 11240 30490 11296 30492
rect 10920 30438 10922 30490
rect 10922 30438 10974 30490
rect 10974 30438 10976 30490
rect 11000 30438 11038 30490
rect 11038 30438 11050 30490
rect 11050 30438 11056 30490
rect 11080 30438 11102 30490
rect 11102 30438 11114 30490
rect 11114 30438 11136 30490
rect 11160 30438 11166 30490
rect 11166 30438 11178 30490
rect 11178 30438 11216 30490
rect 11240 30438 11242 30490
rect 11242 30438 11294 30490
rect 11294 30438 11296 30490
rect 10920 30436 10976 30438
rect 11000 30436 11056 30438
rect 11080 30436 11136 30438
rect 11160 30436 11216 30438
rect 11240 30436 11296 30438
rect 10180 29946 10236 29948
rect 10260 29946 10316 29948
rect 10340 29946 10396 29948
rect 10420 29946 10476 29948
rect 10500 29946 10556 29948
rect 10180 29894 10182 29946
rect 10182 29894 10234 29946
rect 10234 29894 10236 29946
rect 10260 29894 10298 29946
rect 10298 29894 10310 29946
rect 10310 29894 10316 29946
rect 10340 29894 10362 29946
rect 10362 29894 10374 29946
rect 10374 29894 10396 29946
rect 10420 29894 10426 29946
rect 10426 29894 10438 29946
rect 10438 29894 10476 29946
rect 10500 29894 10502 29946
rect 10502 29894 10554 29946
rect 10554 29894 10556 29946
rect 10180 29892 10236 29894
rect 10260 29892 10316 29894
rect 10340 29892 10396 29894
rect 10420 29892 10476 29894
rect 10500 29892 10556 29894
rect 10180 28858 10236 28860
rect 10260 28858 10316 28860
rect 10340 28858 10396 28860
rect 10420 28858 10476 28860
rect 10500 28858 10556 28860
rect 10180 28806 10182 28858
rect 10182 28806 10234 28858
rect 10234 28806 10236 28858
rect 10260 28806 10298 28858
rect 10298 28806 10310 28858
rect 10310 28806 10316 28858
rect 10340 28806 10362 28858
rect 10362 28806 10374 28858
rect 10374 28806 10396 28858
rect 10420 28806 10426 28858
rect 10426 28806 10438 28858
rect 10438 28806 10476 28858
rect 10500 28806 10502 28858
rect 10502 28806 10554 28858
rect 10554 28806 10556 28858
rect 10180 28804 10236 28806
rect 10260 28804 10316 28806
rect 10340 28804 10396 28806
rect 10420 28804 10476 28806
rect 10500 28804 10556 28806
rect 10180 27770 10236 27772
rect 10260 27770 10316 27772
rect 10340 27770 10396 27772
rect 10420 27770 10476 27772
rect 10500 27770 10556 27772
rect 10180 27718 10182 27770
rect 10182 27718 10234 27770
rect 10234 27718 10236 27770
rect 10260 27718 10298 27770
rect 10298 27718 10310 27770
rect 10310 27718 10316 27770
rect 10340 27718 10362 27770
rect 10362 27718 10374 27770
rect 10374 27718 10396 27770
rect 10420 27718 10426 27770
rect 10426 27718 10438 27770
rect 10438 27718 10476 27770
rect 10500 27718 10502 27770
rect 10502 27718 10554 27770
rect 10554 27718 10556 27770
rect 10180 27716 10236 27718
rect 10260 27716 10316 27718
rect 10340 27716 10396 27718
rect 10420 27716 10476 27718
rect 10500 27716 10556 27718
rect 10180 26682 10236 26684
rect 10260 26682 10316 26684
rect 10340 26682 10396 26684
rect 10420 26682 10476 26684
rect 10500 26682 10556 26684
rect 10180 26630 10182 26682
rect 10182 26630 10234 26682
rect 10234 26630 10236 26682
rect 10260 26630 10298 26682
rect 10298 26630 10310 26682
rect 10310 26630 10316 26682
rect 10340 26630 10362 26682
rect 10362 26630 10374 26682
rect 10374 26630 10396 26682
rect 10420 26630 10426 26682
rect 10426 26630 10438 26682
rect 10438 26630 10476 26682
rect 10500 26630 10502 26682
rect 10502 26630 10554 26682
rect 10554 26630 10556 26682
rect 10180 26628 10236 26630
rect 10260 26628 10316 26630
rect 10340 26628 10396 26630
rect 10420 26628 10476 26630
rect 10500 26628 10556 26630
rect 10920 29402 10976 29404
rect 11000 29402 11056 29404
rect 11080 29402 11136 29404
rect 11160 29402 11216 29404
rect 11240 29402 11296 29404
rect 10920 29350 10922 29402
rect 10922 29350 10974 29402
rect 10974 29350 10976 29402
rect 11000 29350 11038 29402
rect 11038 29350 11050 29402
rect 11050 29350 11056 29402
rect 11080 29350 11102 29402
rect 11102 29350 11114 29402
rect 11114 29350 11136 29402
rect 11160 29350 11166 29402
rect 11166 29350 11178 29402
rect 11178 29350 11216 29402
rect 11240 29350 11242 29402
rect 11242 29350 11294 29402
rect 11294 29350 11296 29402
rect 10920 29348 10976 29350
rect 11000 29348 11056 29350
rect 11080 29348 11136 29350
rect 11160 29348 11216 29350
rect 11240 29348 11296 29350
rect 10920 28314 10976 28316
rect 11000 28314 11056 28316
rect 11080 28314 11136 28316
rect 11160 28314 11216 28316
rect 11240 28314 11296 28316
rect 10920 28262 10922 28314
rect 10922 28262 10974 28314
rect 10974 28262 10976 28314
rect 11000 28262 11038 28314
rect 11038 28262 11050 28314
rect 11050 28262 11056 28314
rect 11080 28262 11102 28314
rect 11102 28262 11114 28314
rect 11114 28262 11136 28314
rect 11160 28262 11166 28314
rect 11166 28262 11178 28314
rect 11178 28262 11216 28314
rect 11240 28262 11242 28314
rect 11242 28262 11294 28314
rect 11294 28262 11296 28314
rect 10920 28260 10976 28262
rect 11000 28260 11056 28262
rect 11080 28260 11136 28262
rect 11160 28260 11216 28262
rect 11240 28260 11296 28262
rect 16180 31034 16236 31036
rect 16260 31034 16316 31036
rect 16340 31034 16396 31036
rect 16420 31034 16476 31036
rect 16500 31034 16556 31036
rect 16180 30982 16182 31034
rect 16182 30982 16234 31034
rect 16234 30982 16236 31034
rect 16260 30982 16298 31034
rect 16298 30982 16310 31034
rect 16310 30982 16316 31034
rect 16340 30982 16362 31034
rect 16362 30982 16374 31034
rect 16374 30982 16396 31034
rect 16420 30982 16426 31034
rect 16426 30982 16438 31034
rect 16438 30982 16476 31034
rect 16500 30982 16502 31034
rect 16502 30982 16554 31034
rect 16554 30982 16556 31034
rect 16180 30980 16236 30982
rect 16260 30980 16316 30982
rect 16340 30980 16396 30982
rect 16420 30980 16476 30982
rect 16500 30980 16556 30982
rect 10920 27226 10976 27228
rect 11000 27226 11056 27228
rect 11080 27226 11136 27228
rect 11160 27226 11216 27228
rect 11240 27226 11296 27228
rect 10920 27174 10922 27226
rect 10922 27174 10974 27226
rect 10974 27174 10976 27226
rect 11000 27174 11038 27226
rect 11038 27174 11050 27226
rect 11050 27174 11056 27226
rect 11080 27174 11102 27226
rect 11102 27174 11114 27226
rect 11114 27174 11136 27226
rect 11160 27174 11166 27226
rect 11166 27174 11178 27226
rect 11178 27174 11216 27226
rect 11240 27174 11242 27226
rect 11242 27174 11294 27226
rect 11294 27174 11296 27226
rect 10920 27172 10976 27174
rect 11000 27172 11056 27174
rect 11080 27172 11136 27174
rect 11160 27172 11216 27174
rect 11240 27172 11296 27174
rect 10920 26138 10976 26140
rect 11000 26138 11056 26140
rect 11080 26138 11136 26140
rect 11160 26138 11216 26140
rect 11240 26138 11296 26140
rect 10920 26086 10922 26138
rect 10922 26086 10974 26138
rect 10974 26086 10976 26138
rect 11000 26086 11038 26138
rect 11038 26086 11050 26138
rect 11050 26086 11056 26138
rect 11080 26086 11102 26138
rect 11102 26086 11114 26138
rect 11114 26086 11136 26138
rect 11160 26086 11166 26138
rect 11166 26086 11178 26138
rect 11178 26086 11216 26138
rect 11240 26086 11242 26138
rect 11242 26086 11294 26138
rect 11294 26086 11296 26138
rect 10920 26084 10976 26086
rect 11000 26084 11056 26086
rect 11080 26084 11136 26086
rect 11160 26084 11216 26086
rect 11240 26084 11296 26086
rect 10180 25594 10236 25596
rect 10260 25594 10316 25596
rect 10340 25594 10396 25596
rect 10420 25594 10476 25596
rect 10500 25594 10556 25596
rect 10180 25542 10182 25594
rect 10182 25542 10234 25594
rect 10234 25542 10236 25594
rect 10260 25542 10298 25594
rect 10298 25542 10310 25594
rect 10310 25542 10316 25594
rect 10340 25542 10362 25594
rect 10362 25542 10374 25594
rect 10374 25542 10396 25594
rect 10420 25542 10426 25594
rect 10426 25542 10438 25594
rect 10438 25542 10476 25594
rect 10500 25542 10502 25594
rect 10502 25542 10554 25594
rect 10554 25542 10556 25594
rect 10180 25540 10236 25542
rect 10260 25540 10316 25542
rect 10340 25540 10396 25542
rect 10420 25540 10476 25542
rect 10500 25540 10556 25542
rect 4180 8186 4236 8188
rect 4260 8186 4316 8188
rect 4340 8186 4396 8188
rect 4420 8186 4476 8188
rect 4500 8186 4556 8188
rect 4180 8134 4182 8186
rect 4182 8134 4234 8186
rect 4234 8134 4236 8186
rect 4260 8134 4298 8186
rect 4298 8134 4310 8186
rect 4310 8134 4316 8186
rect 4340 8134 4362 8186
rect 4362 8134 4374 8186
rect 4374 8134 4396 8186
rect 4420 8134 4426 8186
rect 4426 8134 4438 8186
rect 4438 8134 4476 8186
rect 4500 8134 4502 8186
rect 4502 8134 4554 8186
rect 4554 8134 4556 8186
rect 4180 8132 4236 8134
rect 4260 8132 4316 8134
rect 4340 8132 4396 8134
rect 4420 8132 4476 8134
rect 4500 8132 4556 8134
rect 4920 7642 4976 7644
rect 5000 7642 5056 7644
rect 5080 7642 5136 7644
rect 5160 7642 5216 7644
rect 5240 7642 5296 7644
rect 4920 7590 4922 7642
rect 4922 7590 4974 7642
rect 4974 7590 4976 7642
rect 5000 7590 5038 7642
rect 5038 7590 5050 7642
rect 5050 7590 5056 7642
rect 5080 7590 5102 7642
rect 5102 7590 5114 7642
rect 5114 7590 5136 7642
rect 5160 7590 5166 7642
rect 5166 7590 5178 7642
rect 5178 7590 5216 7642
rect 5240 7590 5242 7642
rect 5242 7590 5294 7642
rect 5294 7590 5296 7642
rect 4920 7588 4976 7590
rect 5000 7588 5056 7590
rect 5080 7588 5136 7590
rect 5160 7588 5216 7590
rect 5240 7588 5296 7590
rect 4180 7098 4236 7100
rect 4260 7098 4316 7100
rect 4340 7098 4396 7100
rect 4420 7098 4476 7100
rect 4500 7098 4556 7100
rect 4180 7046 4182 7098
rect 4182 7046 4234 7098
rect 4234 7046 4236 7098
rect 4260 7046 4298 7098
rect 4298 7046 4310 7098
rect 4310 7046 4316 7098
rect 4340 7046 4362 7098
rect 4362 7046 4374 7098
rect 4374 7046 4396 7098
rect 4420 7046 4426 7098
rect 4426 7046 4438 7098
rect 4438 7046 4476 7098
rect 4500 7046 4502 7098
rect 4502 7046 4554 7098
rect 4554 7046 4556 7098
rect 4180 7044 4236 7046
rect 4260 7044 4316 7046
rect 4340 7044 4396 7046
rect 4420 7044 4476 7046
rect 4500 7044 4556 7046
rect 4920 6554 4976 6556
rect 5000 6554 5056 6556
rect 5080 6554 5136 6556
rect 5160 6554 5216 6556
rect 5240 6554 5296 6556
rect 4920 6502 4922 6554
rect 4922 6502 4974 6554
rect 4974 6502 4976 6554
rect 5000 6502 5038 6554
rect 5038 6502 5050 6554
rect 5050 6502 5056 6554
rect 5080 6502 5102 6554
rect 5102 6502 5114 6554
rect 5114 6502 5136 6554
rect 5160 6502 5166 6554
rect 5166 6502 5178 6554
rect 5178 6502 5216 6554
rect 5240 6502 5242 6554
rect 5242 6502 5294 6554
rect 5294 6502 5296 6554
rect 4920 6500 4976 6502
rect 5000 6500 5056 6502
rect 5080 6500 5136 6502
rect 5160 6500 5216 6502
rect 5240 6500 5296 6502
rect 4180 6010 4236 6012
rect 4260 6010 4316 6012
rect 4340 6010 4396 6012
rect 4420 6010 4476 6012
rect 4500 6010 4556 6012
rect 4180 5958 4182 6010
rect 4182 5958 4234 6010
rect 4234 5958 4236 6010
rect 4260 5958 4298 6010
rect 4298 5958 4310 6010
rect 4310 5958 4316 6010
rect 4340 5958 4362 6010
rect 4362 5958 4374 6010
rect 4374 5958 4396 6010
rect 4420 5958 4426 6010
rect 4426 5958 4438 6010
rect 4438 5958 4476 6010
rect 4500 5958 4502 6010
rect 4502 5958 4554 6010
rect 4554 5958 4556 6010
rect 4180 5956 4236 5958
rect 4260 5956 4316 5958
rect 4340 5956 4396 5958
rect 4420 5956 4476 5958
rect 4500 5956 4556 5958
rect 8022 17040 8078 17096
rect 9678 20984 9734 21040
rect 9586 17584 9642 17640
rect 10180 24506 10236 24508
rect 10260 24506 10316 24508
rect 10340 24506 10396 24508
rect 10420 24506 10476 24508
rect 10500 24506 10556 24508
rect 10180 24454 10182 24506
rect 10182 24454 10234 24506
rect 10234 24454 10236 24506
rect 10260 24454 10298 24506
rect 10298 24454 10310 24506
rect 10310 24454 10316 24506
rect 10340 24454 10362 24506
rect 10362 24454 10374 24506
rect 10374 24454 10396 24506
rect 10420 24454 10426 24506
rect 10426 24454 10438 24506
rect 10438 24454 10476 24506
rect 10500 24454 10502 24506
rect 10502 24454 10554 24506
rect 10554 24454 10556 24506
rect 10180 24452 10236 24454
rect 10260 24452 10316 24454
rect 10340 24452 10396 24454
rect 10420 24452 10476 24454
rect 10500 24452 10556 24454
rect 10920 25050 10976 25052
rect 11000 25050 11056 25052
rect 11080 25050 11136 25052
rect 11160 25050 11216 25052
rect 11240 25050 11296 25052
rect 10920 24998 10922 25050
rect 10922 24998 10974 25050
rect 10974 24998 10976 25050
rect 11000 24998 11038 25050
rect 11038 24998 11050 25050
rect 11050 24998 11056 25050
rect 11080 24998 11102 25050
rect 11102 24998 11114 25050
rect 11114 24998 11136 25050
rect 11160 24998 11166 25050
rect 11166 24998 11178 25050
rect 11178 24998 11216 25050
rect 11240 24998 11242 25050
rect 11242 24998 11294 25050
rect 11294 24998 11296 25050
rect 10920 24996 10976 24998
rect 11000 24996 11056 24998
rect 11080 24996 11136 24998
rect 11160 24996 11216 24998
rect 11240 24996 11296 24998
rect 10690 23568 10746 23624
rect 10920 23962 10976 23964
rect 11000 23962 11056 23964
rect 11080 23962 11136 23964
rect 11160 23962 11216 23964
rect 11240 23962 11296 23964
rect 10920 23910 10922 23962
rect 10922 23910 10974 23962
rect 10974 23910 10976 23962
rect 11000 23910 11038 23962
rect 11038 23910 11050 23962
rect 11050 23910 11056 23962
rect 11080 23910 11102 23962
rect 11102 23910 11114 23962
rect 11114 23910 11136 23962
rect 11160 23910 11166 23962
rect 11166 23910 11178 23962
rect 11178 23910 11216 23962
rect 11240 23910 11242 23962
rect 11242 23910 11294 23962
rect 11294 23910 11296 23962
rect 10920 23908 10976 23910
rect 11000 23908 11056 23910
rect 11080 23908 11136 23910
rect 11160 23908 11216 23910
rect 11240 23908 11296 23910
rect 10180 23418 10236 23420
rect 10260 23418 10316 23420
rect 10340 23418 10396 23420
rect 10420 23418 10476 23420
rect 10500 23418 10556 23420
rect 10180 23366 10182 23418
rect 10182 23366 10234 23418
rect 10234 23366 10236 23418
rect 10260 23366 10298 23418
rect 10298 23366 10310 23418
rect 10310 23366 10316 23418
rect 10340 23366 10362 23418
rect 10362 23366 10374 23418
rect 10374 23366 10396 23418
rect 10420 23366 10426 23418
rect 10426 23366 10438 23418
rect 10438 23366 10476 23418
rect 10500 23366 10502 23418
rect 10502 23366 10554 23418
rect 10554 23366 10556 23418
rect 10180 23364 10236 23366
rect 10260 23364 10316 23366
rect 10340 23364 10396 23366
rect 10420 23364 10476 23366
rect 10500 23364 10556 23366
rect 10230 23060 10232 23080
rect 10232 23060 10284 23080
rect 10284 23060 10286 23080
rect 10230 23024 10286 23060
rect 10180 22330 10236 22332
rect 10260 22330 10316 22332
rect 10340 22330 10396 22332
rect 10420 22330 10476 22332
rect 10500 22330 10556 22332
rect 10180 22278 10182 22330
rect 10182 22278 10234 22330
rect 10234 22278 10236 22330
rect 10260 22278 10298 22330
rect 10298 22278 10310 22330
rect 10310 22278 10316 22330
rect 10340 22278 10362 22330
rect 10362 22278 10374 22330
rect 10374 22278 10396 22330
rect 10420 22278 10426 22330
rect 10426 22278 10438 22330
rect 10438 22278 10476 22330
rect 10500 22278 10502 22330
rect 10502 22278 10554 22330
rect 10554 22278 10556 22330
rect 10180 22276 10236 22278
rect 10260 22276 10316 22278
rect 10340 22276 10396 22278
rect 10420 22276 10476 22278
rect 10500 22276 10556 22278
rect 10180 21242 10236 21244
rect 10260 21242 10316 21244
rect 10340 21242 10396 21244
rect 10420 21242 10476 21244
rect 10500 21242 10556 21244
rect 10180 21190 10182 21242
rect 10182 21190 10234 21242
rect 10234 21190 10236 21242
rect 10260 21190 10298 21242
rect 10298 21190 10310 21242
rect 10310 21190 10316 21242
rect 10340 21190 10362 21242
rect 10362 21190 10374 21242
rect 10374 21190 10396 21242
rect 10420 21190 10426 21242
rect 10426 21190 10438 21242
rect 10438 21190 10476 21242
rect 10500 21190 10502 21242
rect 10502 21190 10554 21242
rect 10554 21190 10556 21242
rect 10180 21188 10236 21190
rect 10260 21188 10316 21190
rect 10340 21188 10396 21190
rect 10420 21188 10476 21190
rect 10500 21188 10556 21190
rect 10322 20984 10378 21040
rect 10920 22874 10976 22876
rect 11000 22874 11056 22876
rect 11080 22874 11136 22876
rect 11160 22874 11216 22876
rect 11240 22874 11296 22876
rect 10920 22822 10922 22874
rect 10922 22822 10974 22874
rect 10974 22822 10976 22874
rect 11000 22822 11038 22874
rect 11038 22822 11050 22874
rect 11050 22822 11056 22874
rect 11080 22822 11102 22874
rect 11102 22822 11114 22874
rect 11114 22822 11136 22874
rect 11160 22822 11166 22874
rect 11166 22822 11178 22874
rect 11178 22822 11216 22874
rect 11240 22822 11242 22874
rect 11242 22822 11294 22874
rect 11294 22822 11296 22874
rect 10920 22820 10976 22822
rect 11000 22820 11056 22822
rect 11080 22820 11136 22822
rect 11160 22820 11216 22822
rect 11240 22820 11296 22822
rect 10598 20848 10654 20904
rect 10180 20154 10236 20156
rect 10260 20154 10316 20156
rect 10340 20154 10396 20156
rect 10420 20154 10476 20156
rect 10500 20154 10556 20156
rect 10180 20102 10182 20154
rect 10182 20102 10234 20154
rect 10234 20102 10236 20154
rect 10260 20102 10298 20154
rect 10298 20102 10310 20154
rect 10310 20102 10316 20154
rect 10340 20102 10362 20154
rect 10362 20102 10374 20154
rect 10374 20102 10396 20154
rect 10420 20102 10426 20154
rect 10426 20102 10438 20154
rect 10438 20102 10476 20154
rect 10500 20102 10502 20154
rect 10502 20102 10554 20154
rect 10554 20102 10556 20154
rect 10180 20100 10236 20102
rect 10260 20100 10316 20102
rect 10340 20100 10396 20102
rect 10420 20100 10476 20102
rect 10500 20100 10556 20102
rect 10920 21786 10976 21788
rect 11000 21786 11056 21788
rect 11080 21786 11136 21788
rect 11160 21786 11216 21788
rect 11240 21786 11296 21788
rect 10920 21734 10922 21786
rect 10922 21734 10974 21786
rect 10974 21734 10976 21786
rect 11000 21734 11038 21786
rect 11038 21734 11050 21786
rect 11050 21734 11056 21786
rect 11080 21734 11102 21786
rect 11102 21734 11114 21786
rect 11114 21734 11136 21786
rect 11160 21734 11166 21786
rect 11166 21734 11178 21786
rect 11178 21734 11216 21786
rect 11240 21734 11242 21786
rect 11242 21734 11294 21786
rect 11294 21734 11296 21786
rect 10920 21732 10976 21734
rect 11000 21732 11056 21734
rect 11080 21732 11136 21734
rect 11160 21732 11216 21734
rect 11240 21732 11296 21734
rect 10920 20698 10976 20700
rect 11000 20698 11056 20700
rect 11080 20698 11136 20700
rect 11160 20698 11216 20700
rect 11240 20698 11296 20700
rect 10920 20646 10922 20698
rect 10922 20646 10974 20698
rect 10974 20646 10976 20698
rect 11000 20646 11038 20698
rect 11038 20646 11050 20698
rect 11050 20646 11056 20698
rect 11080 20646 11102 20698
rect 11102 20646 11114 20698
rect 11114 20646 11136 20698
rect 11160 20646 11166 20698
rect 11166 20646 11178 20698
rect 11178 20646 11216 20698
rect 11240 20646 11242 20698
rect 11242 20646 11294 20698
rect 11294 20646 11296 20698
rect 10920 20644 10976 20646
rect 11000 20644 11056 20646
rect 11080 20644 11136 20646
rect 11160 20644 11216 20646
rect 11240 20644 11296 20646
rect 16920 30490 16976 30492
rect 17000 30490 17056 30492
rect 17080 30490 17136 30492
rect 17160 30490 17216 30492
rect 17240 30490 17296 30492
rect 16920 30438 16922 30490
rect 16922 30438 16974 30490
rect 16974 30438 16976 30490
rect 17000 30438 17038 30490
rect 17038 30438 17050 30490
rect 17050 30438 17056 30490
rect 17080 30438 17102 30490
rect 17102 30438 17114 30490
rect 17114 30438 17136 30490
rect 17160 30438 17166 30490
rect 17166 30438 17178 30490
rect 17178 30438 17216 30490
rect 17240 30438 17242 30490
rect 17242 30438 17294 30490
rect 17294 30438 17296 30490
rect 16920 30436 16976 30438
rect 17000 30436 17056 30438
rect 17080 30436 17136 30438
rect 17160 30436 17216 30438
rect 17240 30436 17296 30438
rect 16180 29946 16236 29948
rect 16260 29946 16316 29948
rect 16340 29946 16396 29948
rect 16420 29946 16476 29948
rect 16500 29946 16556 29948
rect 16180 29894 16182 29946
rect 16182 29894 16234 29946
rect 16234 29894 16236 29946
rect 16260 29894 16298 29946
rect 16298 29894 16310 29946
rect 16310 29894 16316 29946
rect 16340 29894 16362 29946
rect 16362 29894 16374 29946
rect 16374 29894 16396 29946
rect 16420 29894 16426 29946
rect 16426 29894 16438 29946
rect 16438 29894 16476 29946
rect 16500 29894 16502 29946
rect 16502 29894 16554 29946
rect 16554 29894 16556 29946
rect 16180 29892 16236 29894
rect 16260 29892 16316 29894
rect 16340 29892 16396 29894
rect 16420 29892 16476 29894
rect 16500 29892 16556 29894
rect 12622 23060 12624 23080
rect 12624 23060 12676 23080
rect 12676 23060 12678 23080
rect 12622 23024 12678 23060
rect 10920 19610 10976 19612
rect 11000 19610 11056 19612
rect 11080 19610 11136 19612
rect 11160 19610 11216 19612
rect 11240 19610 11296 19612
rect 10920 19558 10922 19610
rect 10922 19558 10974 19610
rect 10974 19558 10976 19610
rect 11000 19558 11038 19610
rect 11038 19558 11050 19610
rect 11050 19558 11056 19610
rect 11080 19558 11102 19610
rect 11102 19558 11114 19610
rect 11114 19558 11136 19610
rect 11160 19558 11166 19610
rect 11166 19558 11178 19610
rect 11178 19558 11216 19610
rect 11240 19558 11242 19610
rect 11242 19558 11294 19610
rect 11294 19558 11296 19610
rect 10920 19556 10976 19558
rect 11000 19556 11056 19558
rect 11080 19556 11136 19558
rect 11160 19556 11216 19558
rect 11240 19556 11296 19558
rect 10180 19066 10236 19068
rect 10260 19066 10316 19068
rect 10340 19066 10396 19068
rect 10420 19066 10476 19068
rect 10500 19066 10556 19068
rect 10180 19014 10182 19066
rect 10182 19014 10234 19066
rect 10234 19014 10236 19066
rect 10260 19014 10298 19066
rect 10298 19014 10310 19066
rect 10310 19014 10316 19066
rect 10340 19014 10362 19066
rect 10362 19014 10374 19066
rect 10374 19014 10396 19066
rect 10420 19014 10426 19066
rect 10426 19014 10438 19066
rect 10438 19014 10476 19066
rect 10500 19014 10502 19066
rect 10502 19014 10554 19066
rect 10554 19014 10556 19066
rect 10180 19012 10236 19014
rect 10260 19012 10316 19014
rect 10340 19012 10396 19014
rect 10420 19012 10476 19014
rect 10500 19012 10556 19014
rect 10920 18522 10976 18524
rect 11000 18522 11056 18524
rect 11080 18522 11136 18524
rect 11160 18522 11216 18524
rect 11240 18522 11296 18524
rect 10920 18470 10922 18522
rect 10922 18470 10974 18522
rect 10974 18470 10976 18522
rect 11000 18470 11038 18522
rect 11038 18470 11050 18522
rect 11050 18470 11056 18522
rect 11080 18470 11102 18522
rect 11102 18470 11114 18522
rect 11114 18470 11136 18522
rect 11160 18470 11166 18522
rect 11166 18470 11178 18522
rect 11178 18470 11216 18522
rect 11240 18470 11242 18522
rect 11242 18470 11294 18522
rect 11294 18470 11296 18522
rect 10920 18468 10976 18470
rect 11000 18468 11056 18470
rect 11080 18468 11136 18470
rect 11160 18468 11216 18470
rect 11240 18468 11296 18470
rect 10180 17978 10236 17980
rect 10260 17978 10316 17980
rect 10340 17978 10396 17980
rect 10420 17978 10476 17980
rect 10500 17978 10556 17980
rect 10180 17926 10182 17978
rect 10182 17926 10234 17978
rect 10234 17926 10236 17978
rect 10260 17926 10298 17978
rect 10298 17926 10310 17978
rect 10310 17926 10316 17978
rect 10340 17926 10362 17978
rect 10362 17926 10374 17978
rect 10374 17926 10396 17978
rect 10420 17926 10426 17978
rect 10426 17926 10438 17978
rect 10438 17926 10476 17978
rect 10500 17926 10502 17978
rect 10502 17926 10554 17978
rect 10554 17926 10556 17978
rect 10180 17924 10236 17926
rect 10260 17924 10316 17926
rect 10340 17924 10396 17926
rect 10420 17924 10476 17926
rect 10500 17924 10556 17926
rect 10920 17434 10976 17436
rect 11000 17434 11056 17436
rect 11080 17434 11136 17436
rect 11160 17434 11216 17436
rect 11240 17434 11296 17436
rect 10920 17382 10922 17434
rect 10922 17382 10974 17434
rect 10974 17382 10976 17434
rect 11000 17382 11038 17434
rect 11038 17382 11050 17434
rect 11050 17382 11056 17434
rect 11080 17382 11102 17434
rect 11102 17382 11114 17434
rect 11114 17382 11136 17434
rect 11160 17382 11166 17434
rect 11166 17382 11178 17434
rect 11178 17382 11216 17434
rect 11240 17382 11242 17434
rect 11242 17382 11294 17434
rect 11294 17382 11296 17434
rect 10920 17380 10976 17382
rect 11000 17380 11056 17382
rect 11080 17380 11136 17382
rect 11160 17380 11216 17382
rect 11240 17380 11296 17382
rect 10180 16890 10236 16892
rect 10260 16890 10316 16892
rect 10340 16890 10396 16892
rect 10420 16890 10476 16892
rect 10500 16890 10556 16892
rect 10180 16838 10182 16890
rect 10182 16838 10234 16890
rect 10234 16838 10236 16890
rect 10260 16838 10298 16890
rect 10298 16838 10310 16890
rect 10310 16838 10316 16890
rect 10340 16838 10362 16890
rect 10362 16838 10374 16890
rect 10374 16838 10396 16890
rect 10420 16838 10426 16890
rect 10426 16838 10438 16890
rect 10438 16838 10476 16890
rect 10500 16838 10502 16890
rect 10502 16838 10554 16890
rect 10554 16838 10556 16890
rect 10180 16836 10236 16838
rect 10260 16836 10316 16838
rect 10340 16836 10396 16838
rect 10420 16836 10476 16838
rect 10500 16836 10556 16838
rect 10874 17176 10930 17232
rect 10180 15802 10236 15804
rect 10260 15802 10316 15804
rect 10340 15802 10396 15804
rect 10420 15802 10476 15804
rect 10500 15802 10556 15804
rect 10180 15750 10182 15802
rect 10182 15750 10234 15802
rect 10234 15750 10236 15802
rect 10260 15750 10298 15802
rect 10298 15750 10310 15802
rect 10310 15750 10316 15802
rect 10340 15750 10362 15802
rect 10362 15750 10374 15802
rect 10374 15750 10396 15802
rect 10420 15750 10426 15802
rect 10426 15750 10438 15802
rect 10438 15750 10476 15802
rect 10500 15750 10502 15802
rect 10502 15750 10554 15802
rect 10554 15750 10556 15802
rect 10180 15748 10236 15750
rect 10260 15748 10316 15750
rect 10340 15748 10396 15750
rect 10420 15748 10476 15750
rect 10500 15748 10556 15750
rect 11426 17312 11482 17368
rect 10920 16346 10976 16348
rect 11000 16346 11056 16348
rect 11080 16346 11136 16348
rect 11160 16346 11216 16348
rect 11240 16346 11296 16348
rect 10920 16294 10922 16346
rect 10922 16294 10974 16346
rect 10974 16294 10976 16346
rect 11000 16294 11038 16346
rect 11038 16294 11050 16346
rect 11050 16294 11056 16346
rect 11080 16294 11102 16346
rect 11102 16294 11114 16346
rect 11114 16294 11136 16346
rect 11160 16294 11166 16346
rect 11166 16294 11178 16346
rect 11178 16294 11216 16346
rect 11240 16294 11242 16346
rect 11242 16294 11294 16346
rect 11294 16294 11296 16346
rect 10920 16292 10976 16294
rect 11000 16292 11056 16294
rect 11080 16292 11136 16294
rect 11160 16292 11216 16294
rect 11240 16292 11296 16294
rect 10180 14714 10236 14716
rect 10260 14714 10316 14716
rect 10340 14714 10396 14716
rect 10420 14714 10476 14716
rect 10500 14714 10556 14716
rect 10180 14662 10182 14714
rect 10182 14662 10234 14714
rect 10234 14662 10236 14714
rect 10260 14662 10298 14714
rect 10298 14662 10310 14714
rect 10310 14662 10316 14714
rect 10340 14662 10362 14714
rect 10362 14662 10374 14714
rect 10374 14662 10396 14714
rect 10420 14662 10426 14714
rect 10426 14662 10438 14714
rect 10438 14662 10476 14714
rect 10500 14662 10502 14714
rect 10502 14662 10554 14714
rect 10554 14662 10556 14714
rect 10180 14660 10236 14662
rect 10260 14660 10316 14662
rect 10340 14660 10396 14662
rect 10420 14660 10476 14662
rect 10500 14660 10556 14662
rect 10180 13626 10236 13628
rect 10260 13626 10316 13628
rect 10340 13626 10396 13628
rect 10420 13626 10476 13628
rect 10500 13626 10556 13628
rect 10180 13574 10182 13626
rect 10182 13574 10234 13626
rect 10234 13574 10236 13626
rect 10260 13574 10298 13626
rect 10298 13574 10310 13626
rect 10310 13574 10316 13626
rect 10340 13574 10362 13626
rect 10362 13574 10374 13626
rect 10374 13574 10396 13626
rect 10420 13574 10426 13626
rect 10426 13574 10438 13626
rect 10438 13574 10476 13626
rect 10500 13574 10502 13626
rect 10502 13574 10554 13626
rect 10554 13574 10556 13626
rect 10180 13572 10236 13574
rect 10260 13572 10316 13574
rect 10340 13572 10396 13574
rect 10420 13572 10476 13574
rect 10500 13572 10556 13574
rect 1398 5480 1454 5536
rect 4920 5466 4976 5468
rect 5000 5466 5056 5468
rect 5080 5466 5136 5468
rect 5160 5466 5216 5468
rect 5240 5466 5296 5468
rect 4920 5414 4922 5466
rect 4922 5414 4974 5466
rect 4974 5414 4976 5466
rect 5000 5414 5038 5466
rect 5038 5414 5050 5466
rect 5050 5414 5056 5466
rect 5080 5414 5102 5466
rect 5102 5414 5114 5466
rect 5114 5414 5136 5466
rect 5160 5414 5166 5466
rect 5166 5414 5178 5466
rect 5178 5414 5216 5466
rect 5240 5414 5242 5466
rect 5242 5414 5294 5466
rect 5294 5414 5296 5466
rect 4920 5412 4976 5414
rect 5000 5412 5056 5414
rect 5080 5412 5136 5414
rect 5160 5412 5216 5414
rect 5240 5412 5296 5414
rect 10506 12844 10562 12880
rect 10506 12824 10508 12844
rect 10508 12824 10560 12844
rect 10560 12824 10562 12844
rect 10180 12538 10236 12540
rect 10260 12538 10316 12540
rect 10340 12538 10396 12540
rect 10420 12538 10476 12540
rect 10500 12538 10556 12540
rect 10180 12486 10182 12538
rect 10182 12486 10234 12538
rect 10234 12486 10236 12538
rect 10260 12486 10298 12538
rect 10298 12486 10310 12538
rect 10310 12486 10316 12538
rect 10340 12486 10362 12538
rect 10362 12486 10374 12538
rect 10374 12486 10396 12538
rect 10420 12486 10426 12538
rect 10426 12486 10438 12538
rect 10438 12486 10476 12538
rect 10500 12486 10502 12538
rect 10502 12486 10554 12538
rect 10554 12486 10556 12538
rect 10180 12484 10236 12486
rect 10260 12484 10316 12486
rect 10340 12484 10396 12486
rect 10420 12484 10476 12486
rect 10500 12484 10556 12486
rect 10920 15258 10976 15260
rect 11000 15258 11056 15260
rect 11080 15258 11136 15260
rect 11160 15258 11216 15260
rect 11240 15258 11296 15260
rect 10920 15206 10922 15258
rect 10922 15206 10974 15258
rect 10974 15206 10976 15258
rect 11000 15206 11038 15258
rect 11038 15206 11050 15258
rect 11050 15206 11056 15258
rect 11080 15206 11102 15258
rect 11102 15206 11114 15258
rect 11114 15206 11136 15258
rect 11160 15206 11166 15258
rect 11166 15206 11178 15258
rect 11178 15206 11216 15258
rect 11240 15206 11242 15258
rect 11242 15206 11294 15258
rect 11294 15206 11296 15258
rect 10920 15204 10976 15206
rect 11000 15204 11056 15206
rect 11080 15204 11136 15206
rect 11160 15204 11216 15206
rect 11240 15204 11296 15206
rect 10920 14170 10976 14172
rect 11000 14170 11056 14172
rect 11080 14170 11136 14172
rect 11160 14170 11216 14172
rect 11240 14170 11296 14172
rect 10920 14118 10922 14170
rect 10922 14118 10974 14170
rect 10974 14118 10976 14170
rect 11000 14118 11038 14170
rect 11038 14118 11050 14170
rect 11050 14118 11056 14170
rect 11080 14118 11102 14170
rect 11102 14118 11114 14170
rect 11114 14118 11136 14170
rect 11160 14118 11166 14170
rect 11166 14118 11178 14170
rect 11178 14118 11216 14170
rect 11240 14118 11242 14170
rect 11242 14118 11294 14170
rect 11294 14118 11296 14170
rect 10920 14116 10976 14118
rect 11000 14116 11056 14118
rect 11080 14116 11136 14118
rect 11160 14116 11216 14118
rect 11240 14116 11296 14118
rect 10920 13082 10976 13084
rect 11000 13082 11056 13084
rect 11080 13082 11136 13084
rect 11160 13082 11216 13084
rect 11240 13082 11296 13084
rect 10920 13030 10922 13082
rect 10922 13030 10974 13082
rect 10974 13030 10976 13082
rect 11000 13030 11038 13082
rect 11038 13030 11050 13082
rect 11050 13030 11056 13082
rect 11080 13030 11102 13082
rect 11102 13030 11114 13082
rect 11114 13030 11136 13082
rect 11160 13030 11166 13082
rect 11166 13030 11178 13082
rect 11178 13030 11216 13082
rect 11240 13030 11242 13082
rect 11242 13030 11294 13082
rect 11294 13030 11296 13082
rect 10920 13028 10976 13030
rect 11000 13028 11056 13030
rect 11080 13028 11136 13030
rect 11160 13028 11216 13030
rect 11240 13028 11296 13030
rect 10180 11450 10236 11452
rect 10260 11450 10316 11452
rect 10340 11450 10396 11452
rect 10420 11450 10476 11452
rect 10500 11450 10556 11452
rect 10180 11398 10182 11450
rect 10182 11398 10234 11450
rect 10234 11398 10236 11450
rect 10260 11398 10298 11450
rect 10298 11398 10310 11450
rect 10310 11398 10316 11450
rect 10340 11398 10362 11450
rect 10362 11398 10374 11450
rect 10374 11398 10396 11450
rect 10420 11398 10426 11450
rect 10426 11398 10438 11450
rect 10438 11398 10476 11450
rect 10500 11398 10502 11450
rect 10502 11398 10554 11450
rect 10554 11398 10556 11450
rect 10180 11396 10236 11398
rect 10260 11396 10316 11398
rect 10340 11396 10396 11398
rect 10420 11396 10476 11398
rect 10500 11396 10556 11398
rect 10180 10362 10236 10364
rect 10260 10362 10316 10364
rect 10340 10362 10396 10364
rect 10420 10362 10476 10364
rect 10500 10362 10556 10364
rect 10180 10310 10182 10362
rect 10182 10310 10234 10362
rect 10234 10310 10236 10362
rect 10260 10310 10298 10362
rect 10298 10310 10310 10362
rect 10310 10310 10316 10362
rect 10340 10310 10362 10362
rect 10362 10310 10374 10362
rect 10374 10310 10396 10362
rect 10420 10310 10426 10362
rect 10426 10310 10438 10362
rect 10438 10310 10476 10362
rect 10500 10310 10502 10362
rect 10502 10310 10554 10362
rect 10554 10310 10556 10362
rect 10180 10308 10236 10310
rect 10260 10308 10316 10310
rect 10340 10308 10396 10310
rect 10420 10308 10476 10310
rect 10500 10308 10556 10310
rect 4180 4922 4236 4924
rect 4260 4922 4316 4924
rect 4340 4922 4396 4924
rect 4420 4922 4476 4924
rect 4500 4922 4556 4924
rect 4180 4870 4182 4922
rect 4182 4870 4234 4922
rect 4234 4870 4236 4922
rect 4260 4870 4298 4922
rect 4298 4870 4310 4922
rect 4310 4870 4316 4922
rect 4340 4870 4362 4922
rect 4362 4870 4374 4922
rect 4374 4870 4396 4922
rect 4420 4870 4426 4922
rect 4426 4870 4438 4922
rect 4438 4870 4476 4922
rect 4500 4870 4502 4922
rect 4502 4870 4554 4922
rect 4554 4870 4556 4922
rect 4180 4868 4236 4870
rect 4260 4868 4316 4870
rect 4340 4868 4396 4870
rect 4420 4868 4476 4870
rect 4500 4868 4556 4870
rect 4920 4378 4976 4380
rect 5000 4378 5056 4380
rect 5080 4378 5136 4380
rect 5160 4378 5216 4380
rect 5240 4378 5296 4380
rect 4920 4326 4922 4378
rect 4922 4326 4974 4378
rect 4974 4326 4976 4378
rect 5000 4326 5038 4378
rect 5038 4326 5050 4378
rect 5050 4326 5056 4378
rect 5080 4326 5102 4378
rect 5102 4326 5114 4378
rect 5114 4326 5136 4378
rect 5160 4326 5166 4378
rect 5166 4326 5178 4378
rect 5178 4326 5216 4378
rect 5240 4326 5242 4378
rect 5242 4326 5294 4378
rect 5294 4326 5296 4378
rect 4920 4324 4976 4326
rect 5000 4324 5056 4326
rect 5080 4324 5136 4326
rect 5160 4324 5216 4326
rect 5240 4324 5296 4326
rect 4180 3834 4236 3836
rect 4260 3834 4316 3836
rect 4340 3834 4396 3836
rect 4420 3834 4476 3836
rect 4500 3834 4556 3836
rect 4180 3782 4182 3834
rect 4182 3782 4234 3834
rect 4234 3782 4236 3834
rect 4260 3782 4298 3834
rect 4298 3782 4310 3834
rect 4310 3782 4316 3834
rect 4340 3782 4362 3834
rect 4362 3782 4374 3834
rect 4374 3782 4396 3834
rect 4420 3782 4426 3834
rect 4426 3782 4438 3834
rect 4438 3782 4476 3834
rect 4500 3782 4502 3834
rect 4502 3782 4554 3834
rect 4554 3782 4556 3834
rect 4180 3780 4236 3782
rect 4260 3780 4316 3782
rect 4340 3780 4396 3782
rect 4420 3780 4476 3782
rect 4500 3780 4556 3782
rect 4920 3290 4976 3292
rect 5000 3290 5056 3292
rect 5080 3290 5136 3292
rect 5160 3290 5216 3292
rect 5240 3290 5296 3292
rect 4920 3238 4922 3290
rect 4922 3238 4974 3290
rect 4974 3238 4976 3290
rect 5000 3238 5038 3290
rect 5038 3238 5050 3290
rect 5050 3238 5056 3290
rect 5080 3238 5102 3290
rect 5102 3238 5114 3290
rect 5114 3238 5136 3290
rect 5160 3238 5166 3290
rect 5166 3238 5178 3290
rect 5178 3238 5216 3290
rect 5240 3238 5242 3290
rect 5242 3238 5294 3290
rect 5294 3238 5296 3290
rect 4920 3236 4976 3238
rect 5000 3236 5056 3238
rect 5080 3236 5136 3238
rect 5160 3236 5216 3238
rect 5240 3236 5296 3238
rect 4180 2746 4236 2748
rect 4260 2746 4316 2748
rect 4340 2746 4396 2748
rect 4420 2746 4476 2748
rect 4500 2746 4556 2748
rect 4180 2694 4182 2746
rect 4182 2694 4234 2746
rect 4234 2694 4236 2746
rect 4260 2694 4298 2746
rect 4298 2694 4310 2746
rect 4310 2694 4316 2746
rect 4340 2694 4362 2746
rect 4362 2694 4374 2746
rect 4374 2694 4396 2746
rect 4420 2694 4426 2746
rect 4426 2694 4438 2746
rect 4438 2694 4476 2746
rect 4500 2694 4502 2746
rect 4502 2694 4554 2746
rect 4554 2694 4556 2746
rect 4180 2692 4236 2694
rect 4260 2692 4316 2694
rect 4340 2692 4396 2694
rect 4420 2692 4476 2694
rect 4500 2692 4556 2694
rect 10180 9274 10236 9276
rect 10260 9274 10316 9276
rect 10340 9274 10396 9276
rect 10420 9274 10476 9276
rect 10500 9274 10556 9276
rect 10180 9222 10182 9274
rect 10182 9222 10234 9274
rect 10234 9222 10236 9274
rect 10260 9222 10298 9274
rect 10298 9222 10310 9274
rect 10310 9222 10316 9274
rect 10340 9222 10362 9274
rect 10362 9222 10374 9274
rect 10374 9222 10396 9274
rect 10420 9222 10426 9274
rect 10426 9222 10438 9274
rect 10438 9222 10476 9274
rect 10500 9222 10502 9274
rect 10502 9222 10554 9274
rect 10554 9222 10556 9274
rect 10180 9220 10236 9222
rect 10260 9220 10316 9222
rect 10340 9220 10396 9222
rect 10420 9220 10476 9222
rect 10500 9220 10556 9222
rect 10920 11994 10976 11996
rect 11000 11994 11056 11996
rect 11080 11994 11136 11996
rect 11160 11994 11216 11996
rect 11240 11994 11296 11996
rect 10920 11942 10922 11994
rect 10922 11942 10974 11994
rect 10974 11942 10976 11994
rect 11000 11942 11038 11994
rect 11038 11942 11050 11994
rect 11050 11942 11056 11994
rect 11080 11942 11102 11994
rect 11102 11942 11114 11994
rect 11114 11942 11136 11994
rect 11160 11942 11166 11994
rect 11166 11942 11178 11994
rect 11178 11942 11216 11994
rect 11240 11942 11242 11994
rect 11242 11942 11294 11994
rect 11294 11942 11296 11994
rect 10920 11940 10976 11942
rect 11000 11940 11056 11942
rect 11080 11940 11136 11942
rect 11160 11940 11216 11942
rect 11240 11940 11296 11942
rect 10920 10906 10976 10908
rect 11000 10906 11056 10908
rect 11080 10906 11136 10908
rect 11160 10906 11216 10908
rect 11240 10906 11296 10908
rect 10920 10854 10922 10906
rect 10922 10854 10974 10906
rect 10974 10854 10976 10906
rect 11000 10854 11038 10906
rect 11038 10854 11050 10906
rect 11050 10854 11056 10906
rect 11080 10854 11102 10906
rect 11102 10854 11114 10906
rect 11114 10854 11136 10906
rect 11160 10854 11166 10906
rect 11166 10854 11178 10906
rect 11178 10854 11216 10906
rect 11240 10854 11242 10906
rect 11242 10854 11294 10906
rect 11294 10854 11296 10906
rect 10920 10852 10976 10854
rect 11000 10852 11056 10854
rect 11080 10852 11136 10854
rect 11160 10852 11216 10854
rect 11240 10852 11296 10854
rect 10920 9818 10976 9820
rect 11000 9818 11056 9820
rect 11080 9818 11136 9820
rect 11160 9818 11216 9820
rect 11240 9818 11296 9820
rect 10920 9766 10922 9818
rect 10922 9766 10974 9818
rect 10974 9766 10976 9818
rect 11000 9766 11038 9818
rect 11038 9766 11050 9818
rect 11050 9766 11056 9818
rect 11080 9766 11102 9818
rect 11102 9766 11114 9818
rect 11114 9766 11136 9818
rect 11160 9766 11166 9818
rect 11166 9766 11178 9818
rect 11178 9766 11216 9818
rect 11240 9766 11242 9818
rect 11242 9766 11294 9818
rect 11294 9766 11296 9818
rect 10920 9764 10976 9766
rect 11000 9764 11056 9766
rect 11080 9764 11136 9766
rect 11160 9764 11216 9766
rect 11240 9764 11296 9766
rect 10920 8730 10976 8732
rect 11000 8730 11056 8732
rect 11080 8730 11136 8732
rect 11160 8730 11216 8732
rect 11240 8730 11296 8732
rect 10920 8678 10922 8730
rect 10922 8678 10974 8730
rect 10974 8678 10976 8730
rect 11000 8678 11038 8730
rect 11038 8678 11050 8730
rect 11050 8678 11056 8730
rect 11080 8678 11102 8730
rect 11102 8678 11114 8730
rect 11114 8678 11136 8730
rect 11160 8678 11166 8730
rect 11166 8678 11178 8730
rect 11178 8678 11216 8730
rect 11240 8678 11242 8730
rect 11242 8678 11294 8730
rect 11294 8678 11296 8730
rect 10920 8676 10976 8678
rect 11000 8676 11056 8678
rect 11080 8676 11136 8678
rect 11160 8676 11216 8678
rect 11240 8676 11296 8678
rect 10180 8186 10236 8188
rect 10260 8186 10316 8188
rect 10340 8186 10396 8188
rect 10420 8186 10476 8188
rect 10500 8186 10556 8188
rect 10180 8134 10182 8186
rect 10182 8134 10234 8186
rect 10234 8134 10236 8186
rect 10260 8134 10298 8186
rect 10298 8134 10310 8186
rect 10310 8134 10316 8186
rect 10340 8134 10362 8186
rect 10362 8134 10374 8186
rect 10374 8134 10396 8186
rect 10420 8134 10426 8186
rect 10426 8134 10438 8186
rect 10438 8134 10476 8186
rect 10500 8134 10502 8186
rect 10502 8134 10554 8186
rect 10554 8134 10556 8186
rect 10180 8132 10236 8134
rect 10260 8132 10316 8134
rect 10340 8132 10396 8134
rect 10420 8132 10476 8134
rect 10500 8132 10556 8134
rect 10180 7098 10236 7100
rect 10260 7098 10316 7100
rect 10340 7098 10396 7100
rect 10420 7098 10476 7100
rect 10500 7098 10556 7100
rect 10180 7046 10182 7098
rect 10182 7046 10234 7098
rect 10234 7046 10236 7098
rect 10260 7046 10298 7098
rect 10298 7046 10310 7098
rect 10310 7046 10316 7098
rect 10340 7046 10362 7098
rect 10362 7046 10374 7098
rect 10374 7046 10396 7098
rect 10420 7046 10426 7098
rect 10426 7046 10438 7098
rect 10438 7046 10476 7098
rect 10500 7046 10502 7098
rect 10502 7046 10554 7098
rect 10554 7046 10556 7098
rect 10180 7044 10236 7046
rect 10260 7044 10316 7046
rect 10340 7044 10396 7046
rect 10420 7044 10476 7046
rect 10500 7044 10556 7046
rect 10920 7642 10976 7644
rect 11000 7642 11056 7644
rect 11080 7642 11136 7644
rect 11160 7642 11216 7644
rect 11240 7642 11296 7644
rect 10920 7590 10922 7642
rect 10922 7590 10974 7642
rect 10974 7590 10976 7642
rect 11000 7590 11038 7642
rect 11038 7590 11050 7642
rect 11050 7590 11056 7642
rect 11080 7590 11102 7642
rect 11102 7590 11114 7642
rect 11114 7590 11136 7642
rect 11160 7590 11166 7642
rect 11166 7590 11178 7642
rect 11178 7590 11216 7642
rect 11240 7590 11242 7642
rect 11242 7590 11294 7642
rect 11294 7590 11296 7642
rect 10920 7588 10976 7590
rect 11000 7588 11056 7590
rect 11080 7588 11136 7590
rect 11160 7588 11216 7590
rect 11240 7588 11296 7590
rect 10920 6554 10976 6556
rect 11000 6554 11056 6556
rect 11080 6554 11136 6556
rect 11160 6554 11216 6556
rect 11240 6554 11296 6556
rect 10920 6502 10922 6554
rect 10922 6502 10974 6554
rect 10974 6502 10976 6554
rect 11000 6502 11038 6554
rect 11038 6502 11050 6554
rect 11050 6502 11056 6554
rect 11080 6502 11102 6554
rect 11102 6502 11114 6554
rect 11114 6502 11136 6554
rect 11160 6502 11166 6554
rect 11166 6502 11178 6554
rect 11178 6502 11216 6554
rect 11240 6502 11242 6554
rect 11242 6502 11294 6554
rect 11294 6502 11296 6554
rect 10920 6500 10976 6502
rect 11000 6500 11056 6502
rect 11080 6500 11136 6502
rect 11160 6500 11216 6502
rect 11240 6500 11296 6502
rect 10180 6010 10236 6012
rect 10260 6010 10316 6012
rect 10340 6010 10396 6012
rect 10420 6010 10476 6012
rect 10500 6010 10556 6012
rect 10180 5958 10182 6010
rect 10182 5958 10234 6010
rect 10234 5958 10236 6010
rect 10260 5958 10298 6010
rect 10298 5958 10310 6010
rect 10310 5958 10316 6010
rect 10340 5958 10362 6010
rect 10362 5958 10374 6010
rect 10374 5958 10396 6010
rect 10420 5958 10426 6010
rect 10426 5958 10438 6010
rect 10438 5958 10476 6010
rect 10500 5958 10502 6010
rect 10502 5958 10554 6010
rect 10554 5958 10556 6010
rect 10180 5956 10236 5958
rect 10260 5956 10316 5958
rect 10340 5956 10396 5958
rect 10420 5956 10476 5958
rect 10500 5956 10556 5958
rect 10180 4922 10236 4924
rect 10260 4922 10316 4924
rect 10340 4922 10396 4924
rect 10420 4922 10476 4924
rect 10500 4922 10556 4924
rect 10180 4870 10182 4922
rect 10182 4870 10234 4922
rect 10234 4870 10236 4922
rect 10260 4870 10298 4922
rect 10298 4870 10310 4922
rect 10310 4870 10316 4922
rect 10340 4870 10362 4922
rect 10362 4870 10374 4922
rect 10374 4870 10396 4922
rect 10420 4870 10426 4922
rect 10426 4870 10438 4922
rect 10438 4870 10476 4922
rect 10500 4870 10502 4922
rect 10502 4870 10554 4922
rect 10554 4870 10556 4922
rect 10180 4868 10236 4870
rect 10260 4868 10316 4870
rect 10340 4868 10396 4870
rect 10420 4868 10476 4870
rect 10500 4868 10556 4870
rect 16920 29402 16976 29404
rect 17000 29402 17056 29404
rect 17080 29402 17136 29404
rect 17160 29402 17216 29404
rect 17240 29402 17296 29404
rect 16920 29350 16922 29402
rect 16922 29350 16974 29402
rect 16974 29350 16976 29402
rect 17000 29350 17038 29402
rect 17038 29350 17050 29402
rect 17050 29350 17056 29402
rect 17080 29350 17102 29402
rect 17102 29350 17114 29402
rect 17114 29350 17136 29402
rect 17160 29350 17166 29402
rect 17166 29350 17178 29402
rect 17178 29350 17216 29402
rect 17240 29350 17242 29402
rect 17242 29350 17294 29402
rect 17294 29350 17296 29402
rect 16920 29348 16976 29350
rect 17000 29348 17056 29350
rect 17080 29348 17136 29350
rect 17160 29348 17216 29350
rect 17240 29348 17296 29350
rect 16180 28858 16236 28860
rect 16260 28858 16316 28860
rect 16340 28858 16396 28860
rect 16420 28858 16476 28860
rect 16500 28858 16556 28860
rect 16180 28806 16182 28858
rect 16182 28806 16234 28858
rect 16234 28806 16236 28858
rect 16260 28806 16298 28858
rect 16298 28806 16310 28858
rect 16310 28806 16316 28858
rect 16340 28806 16362 28858
rect 16362 28806 16374 28858
rect 16374 28806 16396 28858
rect 16420 28806 16426 28858
rect 16426 28806 16438 28858
rect 16438 28806 16476 28858
rect 16500 28806 16502 28858
rect 16502 28806 16554 28858
rect 16554 28806 16556 28858
rect 16180 28804 16236 28806
rect 16260 28804 16316 28806
rect 16340 28804 16396 28806
rect 16420 28804 16476 28806
rect 16500 28804 16556 28806
rect 14738 18708 14740 18728
rect 14740 18708 14792 18728
rect 14792 18708 14794 18728
rect 12254 17720 12310 17776
rect 13450 17076 13452 17096
rect 13452 17076 13504 17096
rect 13504 17076 13506 17096
rect 13450 17040 13506 17076
rect 14738 18672 14794 18708
rect 14462 17312 14518 17368
rect 15198 17756 15200 17776
rect 15200 17756 15252 17776
rect 15252 17756 15254 17776
rect 15198 17720 15254 17756
rect 15198 17332 15254 17368
rect 15198 17312 15200 17332
rect 15200 17312 15252 17332
rect 15252 17312 15254 17332
rect 14738 17176 14794 17232
rect 10920 5466 10976 5468
rect 11000 5466 11056 5468
rect 11080 5466 11136 5468
rect 11160 5466 11216 5468
rect 11240 5466 11296 5468
rect 10920 5414 10922 5466
rect 10922 5414 10974 5466
rect 10974 5414 10976 5466
rect 11000 5414 11038 5466
rect 11038 5414 11050 5466
rect 11050 5414 11056 5466
rect 11080 5414 11102 5466
rect 11102 5414 11114 5466
rect 11114 5414 11136 5466
rect 11160 5414 11166 5466
rect 11166 5414 11178 5466
rect 11178 5414 11216 5466
rect 11240 5414 11242 5466
rect 11242 5414 11294 5466
rect 11294 5414 11296 5466
rect 10920 5412 10976 5414
rect 11000 5412 11056 5414
rect 11080 5412 11136 5414
rect 11160 5412 11216 5414
rect 11240 5412 11296 5414
rect 10180 3834 10236 3836
rect 10260 3834 10316 3836
rect 10340 3834 10396 3836
rect 10420 3834 10476 3836
rect 10500 3834 10556 3836
rect 10180 3782 10182 3834
rect 10182 3782 10234 3834
rect 10234 3782 10236 3834
rect 10260 3782 10298 3834
rect 10298 3782 10310 3834
rect 10310 3782 10316 3834
rect 10340 3782 10362 3834
rect 10362 3782 10374 3834
rect 10374 3782 10396 3834
rect 10420 3782 10426 3834
rect 10426 3782 10438 3834
rect 10438 3782 10476 3834
rect 10500 3782 10502 3834
rect 10502 3782 10554 3834
rect 10554 3782 10556 3834
rect 10180 3780 10236 3782
rect 10260 3780 10316 3782
rect 10340 3780 10396 3782
rect 10420 3780 10476 3782
rect 10500 3780 10556 3782
rect 10920 4378 10976 4380
rect 11000 4378 11056 4380
rect 11080 4378 11136 4380
rect 11160 4378 11216 4380
rect 11240 4378 11296 4380
rect 10920 4326 10922 4378
rect 10922 4326 10974 4378
rect 10974 4326 10976 4378
rect 11000 4326 11038 4378
rect 11038 4326 11050 4378
rect 11050 4326 11056 4378
rect 11080 4326 11102 4378
rect 11102 4326 11114 4378
rect 11114 4326 11136 4378
rect 11160 4326 11166 4378
rect 11166 4326 11178 4378
rect 11178 4326 11216 4378
rect 11240 4326 11242 4378
rect 11242 4326 11294 4378
rect 11294 4326 11296 4378
rect 10920 4324 10976 4326
rect 11000 4324 11056 4326
rect 11080 4324 11136 4326
rect 11160 4324 11216 4326
rect 11240 4324 11296 4326
rect 10920 3290 10976 3292
rect 11000 3290 11056 3292
rect 11080 3290 11136 3292
rect 11160 3290 11216 3292
rect 11240 3290 11296 3292
rect 10920 3238 10922 3290
rect 10922 3238 10974 3290
rect 10974 3238 10976 3290
rect 11000 3238 11038 3290
rect 11038 3238 11050 3290
rect 11050 3238 11056 3290
rect 11080 3238 11102 3290
rect 11102 3238 11114 3290
rect 11114 3238 11136 3290
rect 11160 3238 11166 3290
rect 11166 3238 11178 3290
rect 11178 3238 11216 3290
rect 11240 3238 11242 3290
rect 11242 3238 11294 3290
rect 11294 3238 11296 3290
rect 10920 3236 10976 3238
rect 11000 3236 11056 3238
rect 11080 3236 11136 3238
rect 11160 3236 11216 3238
rect 11240 3236 11296 3238
rect 10180 2746 10236 2748
rect 10260 2746 10316 2748
rect 10340 2746 10396 2748
rect 10420 2746 10476 2748
rect 10500 2746 10556 2748
rect 10180 2694 10182 2746
rect 10182 2694 10234 2746
rect 10234 2694 10236 2746
rect 10260 2694 10298 2746
rect 10298 2694 10310 2746
rect 10310 2694 10316 2746
rect 10340 2694 10362 2746
rect 10362 2694 10374 2746
rect 10374 2694 10396 2746
rect 10420 2694 10426 2746
rect 10426 2694 10438 2746
rect 10438 2694 10476 2746
rect 10500 2694 10502 2746
rect 10502 2694 10554 2746
rect 10554 2694 10556 2746
rect 10180 2692 10236 2694
rect 10260 2692 10316 2694
rect 10340 2692 10396 2694
rect 10420 2692 10476 2694
rect 10500 2692 10556 2694
rect 16920 28314 16976 28316
rect 17000 28314 17056 28316
rect 17080 28314 17136 28316
rect 17160 28314 17216 28316
rect 17240 28314 17296 28316
rect 16920 28262 16922 28314
rect 16922 28262 16974 28314
rect 16974 28262 16976 28314
rect 17000 28262 17038 28314
rect 17038 28262 17050 28314
rect 17050 28262 17056 28314
rect 17080 28262 17102 28314
rect 17102 28262 17114 28314
rect 17114 28262 17136 28314
rect 17160 28262 17166 28314
rect 17166 28262 17178 28314
rect 17178 28262 17216 28314
rect 17240 28262 17242 28314
rect 17242 28262 17294 28314
rect 17294 28262 17296 28314
rect 16920 28260 16976 28262
rect 17000 28260 17056 28262
rect 17080 28260 17136 28262
rect 17160 28260 17216 28262
rect 17240 28260 17296 28262
rect 16180 27770 16236 27772
rect 16260 27770 16316 27772
rect 16340 27770 16396 27772
rect 16420 27770 16476 27772
rect 16500 27770 16556 27772
rect 16180 27718 16182 27770
rect 16182 27718 16234 27770
rect 16234 27718 16236 27770
rect 16260 27718 16298 27770
rect 16298 27718 16310 27770
rect 16310 27718 16316 27770
rect 16340 27718 16362 27770
rect 16362 27718 16374 27770
rect 16374 27718 16396 27770
rect 16420 27718 16426 27770
rect 16426 27718 16438 27770
rect 16438 27718 16476 27770
rect 16500 27718 16502 27770
rect 16502 27718 16554 27770
rect 16554 27718 16556 27770
rect 16180 27716 16236 27718
rect 16260 27716 16316 27718
rect 16340 27716 16396 27718
rect 16420 27716 16476 27718
rect 16500 27716 16556 27718
rect 16180 26682 16236 26684
rect 16260 26682 16316 26684
rect 16340 26682 16396 26684
rect 16420 26682 16476 26684
rect 16500 26682 16556 26684
rect 16180 26630 16182 26682
rect 16182 26630 16234 26682
rect 16234 26630 16236 26682
rect 16260 26630 16298 26682
rect 16298 26630 16310 26682
rect 16310 26630 16316 26682
rect 16340 26630 16362 26682
rect 16362 26630 16374 26682
rect 16374 26630 16396 26682
rect 16420 26630 16426 26682
rect 16426 26630 16438 26682
rect 16438 26630 16476 26682
rect 16500 26630 16502 26682
rect 16502 26630 16554 26682
rect 16554 26630 16556 26682
rect 16180 26628 16236 26630
rect 16260 26628 16316 26630
rect 16340 26628 16396 26630
rect 16420 26628 16476 26630
rect 16500 26628 16556 26630
rect 16920 27226 16976 27228
rect 17000 27226 17056 27228
rect 17080 27226 17136 27228
rect 17160 27226 17216 27228
rect 17240 27226 17296 27228
rect 16920 27174 16922 27226
rect 16922 27174 16974 27226
rect 16974 27174 16976 27226
rect 17000 27174 17038 27226
rect 17038 27174 17050 27226
rect 17050 27174 17056 27226
rect 17080 27174 17102 27226
rect 17102 27174 17114 27226
rect 17114 27174 17136 27226
rect 17160 27174 17166 27226
rect 17166 27174 17178 27226
rect 17178 27174 17216 27226
rect 17240 27174 17242 27226
rect 17242 27174 17294 27226
rect 17294 27174 17296 27226
rect 16920 27172 16976 27174
rect 17000 27172 17056 27174
rect 17080 27172 17136 27174
rect 17160 27172 17216 27174
rect 17240 27172 17296 27174
rect 16920 26138 16976 26140
rect 17000 26138 17056 26140
rect 17080 26138 17136 26140
rect 17160 26138 17216 26140
rect 17240 26138 17296 26140
rect 16920 26086 16922 26138
rect 16922 26086 16974 26138
rect 16974 26086 16976 26138
rect 17000 26086 17038 26138
rect 17038 26086 17050 26138
rect 17050 26086 17056 26138
rect 17080 26086 17102 26138
rect 17102 26086 17114 26138
rect 17114 26086 17136 26138
rect 17160 26086 17166 26138
rect 17166 26086 17178 26138
rect 17178 26086 17216 26138
rect 17240 26086 17242 26138
rect 17242 26086 17294 26138
rect 17294 26086 17296 26138
rect 16920 26084 16976 26086
rect 17000 26084 17056 26086
rect 17080 26084 17136 26086
rect 17160 26084 17216 26086
rect 17240 26084 17296 26086
rect 16180 25594 16236 25596
rect 16260 25594 16316 25596
rect 16340 25594 16396 25596
rect 16420 25594 16476 25596
rect 16500 25594 16556 25596
rect 16180 25542 16182 25594
rect 16182 25542 16234 25594
rect 16234 25542 16236 25594
rect 16260 25542 16298 25594
rect 16298 25542 16310 25594
rect 16310 25542 16316 25594
rect 16340 25542 16362 25594
rect 16362 25542 16374 25594
rect 16374 25542 16396 25594
rect 16420 25542 16426 25594
rect 16426 25542 16438 25594
rect 16438 25542 16476 25594
rect 16500 25542 16502 25594
rect 16502 25542 16554 25594
rect 16554 25542 16556 25594
rect 16180 25540 16236 25542
rect 16260 25540 16316 25542
rect 16340 25540 16396 25542
rect 16420 25540 16476 25542
rect 16500 25540 16556 25542
rect 16920 25050 16976 25052
rect 17000 25050 17056 25052
rect 17080 25050 17136 25052
rect 17160 25050 17216 25052
rect 17240 25050 17296 25052
rect 16920 24998 16922 25050
rect 16922 24998 16974 25050
rect 16974 24998 16976 25050
rect 17000 24998 17038 25050
rect 17038 24998 17050 25050
rect 17050 24998 17056 25050
rect 17080 24998 17102 25050
rect 17102 24998 17114 25050
rect 17114 24998 17136 25050
rect 17160 24998 17166 25050
rect 17166 24998 17178 25050
rect 17178 24998 17216 25050
rect 17240 24998 17242 25050
rect 17242 24998 17294 25050
rect 17294 24998 17296 25050
rect 16920 24996 16976 24998
rect 17000 24996 17056 24998
rect 17080 24996 17136 24998
rect 17160 24996 17216 24998
rect 17240 24996 17296 24998
rect 16180 24506 16236 24508
rect 16260 24506 16316 24508
rect 16340 24506 16396 24508
rect 16420 24506 16476 24508
rect 16500 24506 16556 24508
rect 16180 24454 16182 24506
rect 16182 24454 16234 24506
rect 16234 24454 16236 24506
rect 16260 24454 16298 24506
rect 16298 24454 16310 24506
rect 16310 24454 16316 24506
rect 16340 24454 16362 24506
rect 16362 24454 16374 24506
rect 16374 24454 16396 24506
rect 16420 24454 16426 24506
rect 16426 24454 16438 24506
rect 16438 24454 16476 24506
rect 16500 24454 16502 24506
rect 16502 24454 16554 24506
rect 16554 24454 16556 24506
rect 16180 24452 16236 24454
rect 16260 24452 16316 24454
rect 16340 24452 16396 24454
rect 16420 24452 16476 24454
rect 16500 24452 16556 24454
rect 16920 23962 16976 23964
rect 17000 23962 17056 23964
rect 17080 23962 17136 23964
rect 17160 23962 17216 23964
rect 17240 23962 17296 23964
rect 16920 23910 16922 23962
rect 16922 23910 16974 23962
rect 16974 23910 16976 23962
rect 17000 23910 17038 23962
rect 17038 23910 17050 23962
rect 17050 23910 17056 23962
rect 17080 23910 17102 23962
rect 17102 23910 17114 23962
rect 17114 23910 17136 23962
rect 17160 23910 17166 23962
rect 17166 23910 17178 23962
rect 17178 23910 17216 23962
rect 17240 23910 17242 23962
rect 17242 23910 17294 23962
rect 17294 23910 17296 23962
rect 16920 23908 16976 23910
rect 17000 23908 17056 23910
rect 17080 23908 17136 23910
rect 17160 23908 17216 23910
rect 17240 23908 17296 23910
rect 17222 23568 17278 23624
rect 16180 23418 16236 23420
rect 16260 23418 16316 23420
rect 16340 23418 16396 23420
rect 16420 23418 16476 23420
rect 16500 23418 16556 23420
rect 16180 23366 16182 23418
rect 16182 23366 16234 23418
rect 16234 23366 16236 23418
rect 16260 23366 16298 23418
rect 16298 23366 16310 23418
rect 16310 23366 16316 23418
rect 16340 23366 16362 23418
rect 16362 23366 16374 23418
rect 16374 23366 16396 23418
rect 16420 23366 16426 23418
rect 16426 23366 16438 23418
rect 16438 23366 16476 23418
rect 16500 23366 16502 23418
rect 16502 23366 16554 23418
rect 16554 23366 16556 23418
rect 16180 23364 16236 23366
rect 16260 23364 16316 23366
rect 16340 23364 16396 23366
rect 16420 23364 16476 23366
rect 16500 23364 16556 23366
rect 17866 23432 17922 23488
rect 16920 22874 16976 22876
rect 17000 22874 17056 22876
rect 17080 22874 17136 22876
rect 17160 22874 17216 22876
rect 17240 22874 17296 22876
rect 16920 22822 16922 22874
rect 16922 22822 16974 22874
rect 16974 22822 16976 22874
rect 17000 22822 17038 22874
rect 17038 22822 17050 22874
rect 17050 22822 17056 22874
rect 17080 22822 17102 22874
rect 17102 22822 17114 22874
rect 17114 22822 17136 22874
rect 17160 22822 17166 22874
rect 17166 22822 17178 22874
rect 17178 22822 17216 22874
rect 17240 22822 17242 22874
rect 17242 22822 17294 22874
rect 17294 22822 17296 22874
rect 16920 22820 16976 22822
rect 17000 22820 17056 22822
rect 17080 22820 17136 22822
rect 17160 22820 17216 22822
rect 17240 22820 17296 22822
rect 16180 22330 16236 22332
rect 16260 22330 16316 22332
rect 16340 22330 16396 22332
rect 16420 22330 16476 22332
rect 16500 22330 16556 22332
rect 16180 22278 16182 22330
rect 16182 22278 16234 22330
rect 16234 22278 16236 22330
rect 16260 22278 16298 22330
rect 16298 22278 16310 22330
rect 16310 22278 16316 22330
rect 16340 22278 16362 22330
rect 16362 22278 16374 22330
rect 16374 22278 16396 22330
rect 16420 22278 16426 22330
rect 16426 22278 16438 22330
rect 16438 22278 16476 22330
rect 16500 22278 16502 22330
rect 16502 22278 16554 22330
rect 16554 22278 16556 22330
rect 16180 22276 16236 22278
rect 16260 22276 16316 22278
rect 16340 22276 16396 22278
rect 16420 22276 16476 22278
rect 16500 22276 16556 22278
rect 16486 21956 16542 21992
rect 16486 21936 16488 21956
rect 16488 21936 16540 21956
rect 16540 21936 16542 21956
rect 16180 21242 16236 21244
rect 16260 21242 16316 21244
rect 16340 21242 16396 21244
rect 16420 21242 16476 21244
rect 16500 21242 16556 21244
rect 16180 21190 16182 21242
rect 16182 21190 16234 21242
rect 16234 21190 16236 21242
rect 16260 21190 16298 21242
rect 16298 21190 16310 21242
rect 16310 21190 16316 21242
rect 16340 21190 16362 21242
rect 16362 21190 16374 21242
rect 16374 21190 16396 21242
rect 16420 21190 16426 21242
rect 16426 21190 16438 21242
rect 16438 21190 16476 21242
rect 16500 21190 16502 21242
rect 16502 21190 16554 21242
rect 16554 21190 16556 21242
rect 16180 21188 16236 21190
rect 16260 21188 16316 21190
rect 16340 21188 16396 21190
rect 16420 21188 16476 21190
rect 16500 21188 16556 21190
rect 17406 21936 17462 21992
rect 16920 21786 16976 21788
rect 17000 21786 17056 21788
rect 17080 21786 17136 21788
rect 17160 21786 17216 21788
rect 17240 21786 17296 21788
rect 16920 21734 16922 21786
rect 16922 21734 16974 21786
rect 16974 21734 16976 21786
rect 17000 21734 17038 21786
rect 17038 21734 17050 21786
rect 17050 21734 17056 21786
rect 17080 21734 17102 21786
rect 17102 21734 17114 21786
rect 17114 21734 17136 21786
rect 17160 21734 17166 21786
rect 17166 21734 17178 21786
rect 17178 21734 17216 21786
rect 17240 21734 17242 21786
rect 17242 21734 17294 21786
rect 17294 21734 17296 21786
rect 16920 21732 16976 21734
rect 17000 21732 17056 21734
rect 17080 21732 17136 21734
rect 17160 21732 17216 21734
rect 17240 21732 17296 21734
rect 15474 19352 15530 19408
rect 16946 20848 17002 20904
rect 16920 20698 16976 20700
rect 17000 20698 17056 20700
rect 17080 20698 17136 20700
rect 17160 20698 17216 20700
rect 17240 20698 17296 20700
rect 16920 20646 16922 20698
rect 16922 20646 16974 20698
rect 16974 20646 16976 20698
rect 17000 20646 17038 20698
rect 17038 20646 17050 20698
rect 17050 20646 17056 20698
rect 17080 20646 17102 20698
rect 17102 20646 17114 20698
rect 17114 20646 17136 20698
rect 17160 20646 17166 20698
rect 17166 20646 17178 20698
rect 17178 20646 17216 20698
rect 17240 20646 17242 20698
rect 17242 20646 17294 20698
rect 17294 20646 17296 20698
rect 16920 20644 16976 20646
rect 17000 20644 17056 20646
rect 17080 20644 17136 20646
rect 17160 20644 17216 20646
rect 17240 20644 17296 20646
rect 15934 19896 15990 19952
rect 16180 20154 16236 20156
rect 16260 20154 16316 20156
rect 16340 20154 16396 20156
rect 16420 20154 16476 20156
rect 16500 20154 16556 20156
rect 16180 20102 16182 20154
rect 16182 20102 16234 20154
rect 16234 20102 16236 20154
rect 16260 20102 16298 20154
rect 16298 20102 16310 20154
rect 16310 20102 16316 20154
rect 16340 20102 16362 20154
rect 16362 20102 16374 20154
rect 16374 20102 16396 20154
rect 16420 20102 16426 20154
rect 16426 20102 16438 20154
rect 16438 20102 16476 20154
rect 16500 20102 16502 20154
rect 16502 20102 16554 20154
rect 16554 20102 16556 20154
rect 16180 20100 16236 20102
rect 16260 20100 16316 20102
rect 16340 20100 16396 20102
rect 16420 20100 16476 20102
rect 16500 20100 16556 20102
rect 16180 19066 16236 19068
rect 16260 19066 16316 19068
rect 16340 19066 16396 19068
rect 16420 19066 16476 19068
rect 16500 19066 16556 19068
rect 16180 19014 16182 19066
rect 16182 19014 16234 19066
rect 16234 19014 16236 19066
rect 16260 19014 16298 19066
rect 16298 19014 16310 19066
rect 16310 19014 16316 19066
rect 16340 19014 16362 19066
rect 16362 19014 16374 19066
rect 16374 19014 16396 19066
rect 16420 19014 16426 19066
rect 16426 19014 16438 19066
rect 16438 19014 16476 19066
rect 16500 19014 16502 19066
rect 16502 19014 16554 19066
rect 16554 19014 16556 19066
rect 16180 19012 16236 19014
rect 16260 19012 16316 19014
rect 16340 19012 16396 19014
rect 16420 19012 16476 19014
rect 16500 19012 16556 19014
rect 16302 18808 16358 18864
rect 15934 17756 15936 17776
rect 15936 17756 15988 17776
rect 15988 17756 15990 17776
rect 15934 17720 15990 17756
rect 15658 17584 15714 17640
rect 16920 19610 16976 19612
rect 17000 19610 17056 19612
rect 17080 19610 17136 19612
rect 17160 19610 17216 19612
rect 17240 19610 17296 19612
rect 16920 19558 16922 19610
rect 16922 19558 16974 19610
rect 16974 19558 16976 19610
rect 17000 19558 17038 19610
rect 17038 19558 17050 19610
rect 17050 19558 17056 19610
rect 17080 19558 17102 19610
rect 17102 19558 17114 19610
rect 17114 19558 17136 19610
rect 17160 19558 17166 19610
rect 17166 19558 17178 19610
rect 17178 19558 17216 19610
rect 17240 19558 17242 19610
rect 17242 19558 17294 19610
rect 17294 19558 17296 19610
rect 16920 19556 16976 19558
rect 17000 19556 17056 19558
rect 17080 19556 17136 19558
rect 17160 19556 17216 19558
rect 17240 19556 17296 19558
rect 16946 19352 17002 19408
rect 16920 18522 16976 18524
rect 17000 18522 17056 18524
rect 17080 18522 17136 18524
rect 17160 18522 17216 18524
rect 17240 18522 17296 18524
rect 16920 18470 16922 18522
rect 16922 18470 16974 18522
rect 16974 18470 16976 18522
rect 17000 18470 17038 18522
rect 17038 18470 17050 18522
rect 17050 18470 17056 18522
rect 17080 18470 17102 18522
rect 17102 18470 17114 18522
rect 17114 18470 17136 18522
rect 17160 18470 17166 18522
rect 17166 18470 17178 18522
rect 17178 18470 17216 18522
rect 17240 18470 17242 18522
rect 17242 18470 17294 18522
rect 17294 18470 17296 18522
rect 16920 18468 16976 18470
rect 17000 18468 17056 18470
rect 17080 18468 17136 18470
rect 17160 18468 17216 18470
rect 17240 18468 17296 18470
rect 16180 17978 16236 17980
rect 16260 17978 16316 17980
rect 16340 17978 16396 17980
rect 16420 17978 16476 17980
rect 16500 17978 16556 17980
rect 16180 17926 16182 17978
rect 16182 17926 16234 17978
rect 16234 17926 16236 17978
rect 16260 17926 16298 17978
rect 16298 17926 16310 17978
rect 16310 17926 16316 17978
rect 16340 17926 16362 17978
rect 16362 17926 16374 17978
rect 16374 17926 16396 17978
rect 16420 17926 16426 17978
rect 16426 17926 16438 17978
rect 16438 17926 16476 17978
rect 16500 17926 16502 17978
rect 16502 17926 16554 17978
rect 16554 17926 16556 17978
rect 16180 17924 16236 17926
rect 16260 17924 16316 17926
rect 16340 17924 16396 17926
rect 16420 17924 16476 17926
rect 16500 17924 16556 17926
rect 16486 17196 16542 17232
rect 16486 17176 16488 17196
rect 16488 17176 16540 17196
rect 16540 17176 16542 17196
rect 17314 17584 17370 17640
rect 16920 17434 16976 17436
rect 17000 17434 17056 17436
rect 17080 17434 17136 17436
rect 17160 17434 17216 17436
rect 17240 17434 17296 17436
rect 16920 17382 16922 17434
rect 16922 17382 16974 17434
rect 16974 17382 16976 17434
rect 17000 17382 17038 17434
rect 17038 17382 17050 17434
rect 17050 17382 17056 17434
rect 17080 17382 17102 17434
rect 17102 17382 17114 17434
rect 17114 17382 17136 17434
rect 17160 17382 17166 17434
rect 17166 17382 17178 17434
rect 17178 17382 17216 17434
rect 17240 17382 17242 17434
rect 17242 17382 17294 17434
rect 17294 17382 17296 17434
rect 16920 17380 16976 17382
rect 17000 17380 17056 17382
rect 17080 17380 17136 17382
rect 17160 17380 17216 17382
rect 17240 17380 17296 17382
rect 16180 16890 16236 16892
rect 16260 16890 16316 16892
rect 16340 16890 16396 16892
rect 16420 16890 16476 16892
rect 16500 16890 16556 16892
rect 16180 16838 16182 16890
rect 16182 16838 16234 16890
rect 16234 16838 16236 16890
rect 16260 16838 16298 16890
rect 16298 16838 16310 16890
rect 16310 16838 16316 16890
rect 16340 16838 16362 16890
rect 16362 16838 16374 16890
rect 16374 16838 16396 16890
rect 16420 16838 16426 16890
rect 16426 16838 16438 16890
rect 16438 16838 16476 16890
rect 16500 16838 16502 16890
rect 16502 16838 16554 16890
rect 16554 16838 16556 16890
rect 16180 16836 16236 16838
rect 16260 16836 16316 16838
rect 16340 16836 16396 16838
rect 16420 16836 16476 16838
rect 16500 16836 16556 16838
rect 16920 16346 16976 16348
rect 17000 16346 17056 16348
rect 17080 16346 17136 16348
rect 17160 16346 17216 16348
rect 17240 16346 17296 16348
rect 16920 16294 16922 16346
rect 16922 16294 16974 16346
rect 16974 16294 16976 16346
rect 17000 16294 17038 16346
rect 17038 16294 17050 16346
rect 17050 16294 17056 16346
rect 17080 16294 17102 16346
rect 17102 16294 17114 16346
rect 17114 16294 17136 16346
rect 17160 16294 17166 16346
rect 17166 16294 17178 16346
rect 17178 16294 17216 16346
rect 17240 16294 17242 16346
rect 17242 16294 17294 16346
rect 17294 16294 17296 16346
rect 16920 16292 16976 16294
rect 17000 16292 17056 16294
rect 17080 16292 17136 16294
rect 17160 16292 17216 16294
rect 17240 16292 17296 16294
rect 15382 11056 15438 11112
rect 16180 15802 16236 15804
rect 16260 15802 16316 15804
rect 16340 15802 16396 15804
rect 16420 15802 16476 15804
rect 16500 15802 16556 15804
rect 16180 15750 16182 15802
rect 16182 15750 16234 15802
rect 16234 15750 16236 15802
rect 16260 15750 16298 15802
rect 16298 15750 16310 15802
rect 16310 15750 16316 15802
rect 16340 15750 16362 15802
rect 16362 15750 16374 15802
rect 16374 15750 16396 15802
rect 16420 15750 16426 15802
rect 16426 15750 16438 15802
rect 16438 15750 16476 15802
rect 16500 15750 16502 15802
rect 16502 15750 16554 15802
rect 16554 15750 16556 15802
rect 16180 15748 16236 15750
rect 16260 15748 16316 15750
rect 16340 15748 16396 15750
rect 16420 15748 16476 15750
rect 16500 15748 16556 15750
rect 16920 15258 16976 15260
rect 17000 15258 17056 15260
rect 17080 15258 17136 15260
rect 17160 15258 17216 15260
rect 17240 15258 17296 15260
rect 16920 15206 16922 15258
rect 16922 15206 16974 15258
rect 16974 15206 16976 15258
rect 17000 15206 17038 15258
rect 17038 15206 17050 15258
rect 17050 15206 17056 15258
rect 17080 15206 17102 15258
rect 17102 15206 17114 15258
rect 17114 15206 17136 15258
rect 17160 15206 17166 15258
rect 17166 15206 17178 15258
rect 17178 15206 17216 15258
rect 17240 15206 17242 15258
rect 17242 15206 17294 15258
rect 17294 15206 17296 15258
rect 16920 15204 16976 15206
rect 17000 15204 17056 15206
rect 17080 15204 17136 15206
rect 17160 15204 17216 15206
rect 17240 15204 17296 15206
rect 16180 14714 16236 14716
rect 16260 14714 16316 14716
rect 16340 14714 16396 14716
rect 16420 14714 16476 14716
rect 16500 14714 16556 14716
rect 16180 14662 16182 14714
rect 16182 14662 16234 14714
rect 16234 14662 16236 14714
rect 16260 14662 16298 14714
rect 16298 14662 16310 14714
rect 16310 14662 16316 14714
rect 16340 14662 16362 14714
rect 16362 14662 16374 14714
rect 16374 14662 16396 14714
rect 16420 14662 16426 14714
rect 16426 14662 16438 14714
rect 16438 14662 16476 14714
rect 16500 14662 16502 14714
rect 16502 14662 16554 14714
rect 16554 14662 16556 14714
rect 16180 14660 16236 14662
rect 16260 14660 16316 14662
rect 16340 14660 16396 14662
rect 16420 14660 16476 14662
rect 16500 14660 16556 14662
rect 16180 13626 16236 13628
rect 16260 13626 16316 13628
rect 16340 13626 16396 13628
rect 16420 13626 16476 13628
rect 16500 13626 16556 13628
rect 16180 13574 16182 13626
rect 16182 13574 16234 13626
rect 16234 13574 16236 13626
rect 16260 13574 16298 13626
rect 16298 13574 16310 13626
rect 16310 13574 16316 13626
rect 16340 13574 16362 13626
rect 16362 13574 16374 13626
rect 16374 13574 16396 13626
rect 16420 13574 16426 13626
rect 16426 13574 16438 13626
rect 16438 13574 16476 13626
rect 16500 13574 16502 13626
rect 16502 13574 16554 13626
rect 16554 13574 16556 13626
rect 16180 13572 16236 13574
rect 16260 13572 16316 13574
rect 16340 13572 16396 13574
rect 16420 13572 16476 13574
rect 16500 13572 16556 13574
rect 16180 12538 16236 12540
rect 16260 12538 16316 12540
rect 16340 12538 16396 12540
rect 16420 12538 16476 12540
rect 16500 12538 16556 12540
rect 16180 12486 16182 12538
rect 16182 12486 16234 12538
rect 16234 12486 16236 12538
rect 16260 12486 16298 12538
rect 16298 12486 16310 12538
rect 16310 12486 16316 12538
rect 16340 12486 16362 12538
rect 16362 12486 16374 12538
rect 16374 12486 16396 12538
rect 16420 12486 16426 12538
rect 16426 12486 16438 12538
rect 16438 12486 16476 12538
rect 16500 12486 16502 12538
rect 16502 12486 16554 12538
rect 16554 12486 16556 12538
rect 16180 12484 16236 12486
rect 16260 12484 16316 12486
rect 16340 12484 16396 12486
rect 16420 12484 16476 12486
rect 16500 12484 16556 12486
rect 16920 14170 16976 14172
rect 17000 14170 17056 14172
rect 17080 14170 17136 14172
rect 17160 14170 17216 14172
rect 17240 14170 17296 14172
rect 16920 14118 16922 14170
rect 16922 14118 16974 14170
rect 16974 14118 16976 14170
rect 17000 14118 17038 14170
rect 17038 14118 17050 14170
rect 17050 14118 17056 14170
rect 17080 14118 17102 14170
rect 17102 14118 17114 14170
rect 17114 14118 17136 14170
rect 17160 14118 17166 14170
rect 17166 14118 17178 14170
rect 17178 14118 17216 14170
rect 17240 14118 17242 14170
rect 17242 14118 17294 14170
rect 17294 14118 17296 14170
rect 16920 14116 16976 14118
rect 17000 14116 17056 14118
rect 17080 14116 17136 14118
rect 17160 14116 17216 14118
rect 17240 14116 17296 14118
rect 16920 13082 16976 13084
rect 17000 13082 17056 13084
rect 17080 13082 17136 13084
rect 17160 13082 17216 13084
rect 17240 13082 17296 13084
rect 16920 13030 16922 13082
rect 16922 13030 16974 13082
rect 16974 13030 16976 13082
rect 17000 13030 17038 13082
rect 17038 13030 17050 13082
rect 17050 13030 17056 13082
rect 17080 13030 17102 13082
rect 17102 13030 17114 13082
rect 17114 13030 17136 13082
rect 17160 13030 17166 13082
rect 17166 13030 17178 13082
rect 17178 13030 17216 13082
rect 17240 13030 17242 13082
rect 17242 13030 17294 13082
rect 17294 13030 17296 13082
rect 16920 13028 16976 13030
rect 17000 13028 17056 13030
rect 17080 13028 17136 13030
rect 17160 13028 17216 13030
rect 17240 13028 17296 13030
rect 17958 18672 18014 18728
rect 16920 11994 16976 11996
rect 17000 11994 17056 11996
rect 17080 11994 17136 11996
rect 17160 11994 17216 11996
rect 17240 11994 17296 11996
rect 16920 11942 16922 11994
rect 16922 11942 16974 11994
rect 16974 11942 16976 11994
rect 17000 11942 17038 11994
rect 17038 11942 17050 11994
rect 17050 11942 17056 11994
rect 17080 11942 17102 11994
rect 17102 11942 17114 11994
rect 17114 11942 17136 11994
rect 17160 11942 17166 11994
rect 17166 11942 17178 11994
rect 17178 11942 17216 11994
rect 17240 11942 17242 11994
rect 17242 11942 17294 11994
rect 17294 11942 17296 11994
rect 16920 11940 16976 11942
rect 17000 11940 17056 11942
rect 17080 11940 17136 11942
rect 17160 11940 17216 11942
rect 17240 11940 17296 11942
rect 16180 11450 16236 11452
rect 16260 11450 16316 11452
rect 16340 11450 16396 11452
rect 16420 11450 16476 11452
rect 16500 11450 16556 11452
rect 16180 11398 16182 11450
rect 16182 11398 16234 11450
rect 16234 11398 16236 11450
rect 16260 11398 16298 11450
rect 16298 11398 16310 11450
rect 16310 11398 16316 11450
rect 16340 11398 16362 11450
rect 16362 11398 16374 11450
rect 16374 11398 16396 11450
rect 16420 11398 16426 11450
rect 16426 11398 16438 11450
rect 16438 11398 16476 11450
rect 16500 11398 16502 11450
rect 16502 11398 16554 11450
rect 16554 11398 16556 11450
rect 16180 11396 16236 11398
rect 16260 11396 16316 11398
rect 16340 11396 16396 11398
rect 16420 11396 16476 11398
rect 16500 11396 16556 11398
rect 16920 10906 16976 10908
rect 17000 10906 17056 10908
rect 17080 10906 17136 10908
rect 17160 10906 17216 10908
rect 17240 10906 17296 10908
rect 16920 10854 16922 10906
rect 16922 10854 16974 10906
rect 16974 10854 16976 10906
rect 17000 10854 17038 10906
rect 17038 10854 17050 10906
rect 17050 10854 17056 10906
rect 17080 10854 17102 10906
rect 17102 10854 17114 10906
rect 17114 10854 17136 10906
rect 17160 10854 17166 10906
rect 17166 10854 17178 10906
rect 17178 10854 17216 10906
rect 17240 10854 17242 10906
rect 17242 10854 17294 10906
rect 17294 10854 17296 10906
rect 16920 10852 16976 10854
rect 17000 10852 17056 10854
rect 17080 10852 17136 10854
rect 17160 10852 17216 10854
rect 17240 10852 17296 10854
rect 16180 10362 16236 10364
rect 16260 10362 16316 10364
rect 16340 10362 16396 10364
rect 16420 10362 16476 10364
rect 16500 10362 16556 10364
rect 16180 10310 16182 10362
rect 16182 10310 16234 10362
rect 16234 10310 16236 10362
rect 16260 10310 16298 10362
rect 16298 10310 16310 10362
rect 16310 10310 16316 10362
rect 16340 10310 16362 10362
rect 16362 10310 16374 10362
rect 16374 10310 16396 10362
rect 16420 10310 16426 10362
rect 16426 10310 16438 10362
rect 16438 10310 16476 10362
rect 16500 10310 16502 10362
rect 16502 10310 16554 10362
rect 16554 10310 16556 10362
rect 16180 10308 16236 10310
rect 16260 10308 16316 10310
rect 16340 10308 16396 10310
rect 16420 10308 16476 10310
rect 16500 10308 16556 10310
rect 16920 9818 16976 9820
rect 17000 9818 17056 9820
rect 17080 9818 17136 9820
rect 17160 9818 17216 9820
rect 17240 9818 17296 9820
rect 16920 9766 16922 9818
rect 16922 9766 16974 9818
rect 16974 9766 16976 9818
rect 17000 9766 17038 9818
rect 17038 9766 17050 9818
rect 17050 9766 17056 9818
rect 17080 9766 17102 9818
rect 17102 9766 17114 9818
rect 17114 9766 17136 9818
rect 17160 9766 17166 9818
rect 17166 9766 17178 9818
rect 17178 9766 17216 9818
rect 17240 9766 17242 9818
rect 17242 9766 17294 9818
rect 17294 9766 17296 9818
rect 16920 9764 16976 9766
rect 17000 9764 17056 9766
rect 17080 9764 17136 9766
rect 17160 9764 17216 9766
rect 17240 9764 17296 9766
rect 16180 9274 16236 9276
rect 16260 9274 16316 9276
rect 16340 9274 16396 9276
rect 16420 9274 16476 9276
rect 16500 9274 16556 9276
rect 16180 9222 16182 9274
rect 16182 9222 16234 9274
rect 16234 9222 16236 9274
rect 16260 9222 16298 9274
rect 16298 9222 16310 9274
rect 16310 9222 16316 9274
rect 16340 9222 16362 9274
rect 16362 9222 16374 9274
rect 16374 9222 16396 9274
rect 16420 9222 16426 9274
rect 16426 9222 16438 9274
rect 16438 9222 16476 9274
rect 16500 9222 16502 9274
rect 16502 9222 16554 9274
rect 16554 9222 16556 9274
rect 16180 9220 16236 9222
rect 16260 9220 16316 9222
rect 16340 9220 16396 9222
rect 16420 9220 16476 9222
rect 16500 9220 16556 9222
rect 16920 8730 16976 8732
rect 17000 8730 17056 8732
rect 17080 8730 17136 8732
rect 17160 8730 17216 8732
rect 17240 8730 17296 8732
rect 16920 8678 16922 8730
rect 16922 8678 16974 8730
rect 16974 8678 16976 8730
rect 17000 8678 17038 8730
rect 17038 8678 17050 8730
rect 17050 8678 17056 8730
rect 17080 8678 17102 8730
rect 17102 8678 17114 8730
rect 17114 8678 17136 8730
rect 17160 8678 17166 8730
rect 17166 8678 17178 8730
rect 17178 8678 17216 8730
rect 17240 8678 17242 8730
rect 17242 8678 17294 8730
rect 17294 8678 17296 8730
rect 16920 8676 16976 8678
rect 17000 8676 17056 8678
rect 17080 8676 17136 8678
rect 17160 8676 17216 8678
rect 17240 8676 17296 8678
rect 16180 8186 16236 8188
rect 16260 8186 16316 8188
rect 16340 8186 16396 8188
rect 16420 8186 16476 8188
rect 16500 8186 16556 8188
rect 16180 8134 16182 8186
rect 16182 8134 16234 8186
rect 16234 8134 16236 8186
rect 16260 8134 16298 8186
rect 16298 8134 16310 8186
rect 16310 8134 16316 8186
rect 16340 8134 16362 8186
rect 16362 8134 16374 8186
rect 16374 8134 16396 8186
rect 16420 8134 16426 8186
rect 16426 8134 16438 8186
rect 16438 8134 16476 8186
rect 16500 8134 16502 8186
rect 16502 8134 16554 8186
rect 16554 8134 16556 8186
rect 16180 8132 16236 8134
rect 16260 8132 16316 8134
rect 16340 8132 16396 8134
rect 16420 8132 16476 8134
rect 16500 8132 16556 8134
rect 24490 31764 24492 31784
rect 24492 31764 24544 31784
rect 24544 31764 24546 31784
rect 24490 31728 24546 31764
rect 22920 31578 22976 31580
rect 23000 31578 23056 31580
rect 23080 31578 23136 31580
rect 23160 31578 23216 31580
rect 23240 31578 23296 31580
rect 22920 31526 22922 31578
rect 22922 31526 22974 31578
rect 22974 31526 22976 31578
rect 23000 31526 23038 31578
rect 23038 31526 23050 31578
rect 23050 31526 23056 31578
rect 23080 31526 23102 31578
rect 23102 31526 23114 31578
rect 23114 31526 23136 31578
rect 23160 31526 23166 31578
rect 23166 31526 23178 31578
rect 23178 31526 23216 31578
rect 23240 31526 23242 31578
rect 23242 31526 23294 31578
rect 23294 31526 23296 31578
rect 22920 31524 22976 31526
rect 23000 31524 23056 31526
rect 23080 31524 23136 31526
rect 23160 31524 23216 31526
rect 23240 31524 23296 31526
rect 18694 26324 18696 26344
rect 18696 26324 18748 26344
rect 18748 26324 18750 26344
rect 18694 26288 18750 26324
rect 19338 23432 19394 23488
rect 19338 20984 19394 21040
rect 18234 18808 18290 18864
rect 19338 19796 19340 19816
rect 19340 19796 19392 19816
rect 19392 19796 19394 19816
rect 19338 19760 19394 19796
rect 20074 19896 20130 19952
rect 19890 19796 19892 19816
rect 19892 19796 19944 19816
rect 19944 19796 19946 19816
rect 19890 19760 19946 19796
rect 22180 31034 22236 31036
rect 22260 31034 22316 31036
rect 22340 31034 22396 31036
rect 22420 31034 22476 31036
rect 22500 31034 22556 31036
rect 22180 30982 22182 31034
rect 22182 30982 22234 31034
rect 22234 30982 22236 31034
rect 22260 30982 22298 31034
rect 22298 30982 22310 31034
rect 22310 30982 22316 31034
rect 22340 30982 22362 31034
rect 22362 30982 22374 31034
rect 22374 30982 22396 31034
rect 22420 30982 22426 31034
rect 22426 30982 22438 31034
rect 22438 30982 22476 31034
rect 22500 30982 22502 31034
rect 22502 30982 22554 31034
rect 22554 30982 22556 31034
rect 22180 30980 22236 30982
rect 22260 30980 22316 30982
rect 22340 30980 22396 30982
rect 22420 30980 22476 30982
rect 22500 30980 22556 30982
rect 22180 29946 22236 29948
rect 22260 29946 22316 29948
rect 22340 29946 22396 29948
rect 22420 29946 22476 29948
rect 22500 29946 22556 29948
rect 22180 29894 22182 29946
rect 22182 29894 22234 29946
rect 22234 29894 22236 29946
rect 22260 29894 22298 29946
rect 22298 29894 22310 29946
rect 22310 29894 22316 29946
rect 22340 29894 22362 29946
rect 22362 29894 22374 29946
rect 22374 29894 22396 29946
rect 22420 29894 22426 29946
rect 22426 29894 22438 29946
rect 22438 29894 22476 29946
rect 22500 29894 22502 29946
rect 22502 29894 22554 29946
rect 22554 29894 22556 29946
rect 22180 29892 22236 29894
rect 22260 29892 22316 29894
rect 22340 29892 22396 29894
rect 22420 29892 22476 29894
rect 22500 29892 22556 29894
rect 22920 30490 22976 30492
rect 23000 30490 23056 30492
rect 23080 30490 23136 30492
rect 23160 30490 23216 30492
rect 23240 30490 23296 30492
rect 22920 30438 22922 30490
rect 22922 30438 22974 30490
rect 22974 30438 22976 30490
rect 23000 30438 23038 30490
rect 23038 30438 23050 30490
rect 23050 30438 23056 30490
rect 23080 30438 23102 30490
rect 23102 30438 23114 30490
rect 23114 30438 23136 30490
rect 23160 30438 23166 30490
rect 23166 30438 23178 30490
rect 23178 30438 23216 30490
rect 23240 30438 23242 30490
rect 23242 30438 23294 30490
rect 23294 30438 23296 30490
rect 22920 30436 22976 30438
rect 23000 30436 23056 30438
rect 23080 30436 23136 30438
rect 23160 30436 23216 30438
rect 23240 30436 23296 30438
rect 22920 29402 22976 29404
rect 23000 29402 23056 29404
rect 23080 29402 23136 29404
rect 23160 29402 23216 29404
rect 23240 29402 23296 29404
rect 22920 29350 22922 29402
rect 22922 29350 22974 29402
rect 22974 29350 22976 29402
rect 23000 29350 23038 29402
rect 23038 29350 23050 29402
rect 23050 29350 23056 29402
rect 23080 29350 23102 29402
rect 23102 29350 23114 29402
rect 23114 29350 23136 29402
rect 23160 29350 23166 29402
rect 23166 29350 23178 29402
rect 23178 29350 23216 29402
rect 23240 29350 23242 29402
rect 23242 29350 23294 29402
rect 23294 29350 23296 29402
rect 22920 29348 22976 29350
rect 23000 29348 23056 29350
rect 23080 29348 23136 29350
rect 23160 29348 23216 29350
rect 23240 29348 23296 29350
rect 22180 28858 22236 28860
rect 22260 28858 22316 28860
rect 22340 28858 22396 28860
rect 22420 28858 22476 28860
rect 22500 28858 22556 28860
rect 22180 28806 22182 28858
rect 22182 28806 22234 28858
rect 22234 28806 22236 28858
rect 22260 28806 22298 28858
rect 22298 28806 22310 28858
rect 22310 28806 22316 28858
rect 22340 28806 22362 28858
rect 22362 28806 22374 28858
rect 22374 28806 22396 28858
rect 22420 28806 22426 28858
rect 22426 28806 22438 28858
rect 22438 28806 22476 28858
rect 22500 28806 22502 28858
rect 22502 28806 22554 28858
rect 22554 28806 22556 28858
rect 22180 28804 22236 28806
rect 22260 28804 22316 28806
rect 22340 28804 22396 28806
rect 22420 28804 22476 28806
rect 22500 28804 22556 28806
rect 22466 27920 22522 27976
rect 22180 27770 22236 27772
rect 22260 27770 22316 27772
rect 22340 27770 22396 27772
rect 22420 27770 22476 27772
rect 22500 27770 22556 27772
rect 22180 27718 22182 27770
rect 22182 27718 22234 27770
rect 22234 27718 22236 27770
rect 22260 27718 22298 27770
rect 22298 27718 22310 27770
rect 22310 27718 22316 27770
rect 22340 27718 22362 27770
rect 22362 27718 22374 27770
rect 22374 27718 22396 27770
rect 22420 27718 22426 27770
rect 22426 27718 22438 27770
rect 22438 27718 22476 27770
rect 22500 27718 22502 27770
rect 22502 27718 22554 27770
rect 22554 27718 22556 27770
rect 22180 27716 22236 27718
rect 22260 27716 22316 27718
rect 22340 27716 22396 27718
rect 22420 27716 22476 27718
rect 22500 27716 22556 27718
rect 22920 28314 22976 28316
rect 23000 28314 23056 28316
rect 23080 28314 23136 28316
rect 23160 28314 23216 28316
rect 23240 28314 23296 28316
rect 22920 28262 22922 28314
rect 22922 28262 22974 28314
rect 22974 28262 22976 28314
rect 23000 28262 23038 28314
rect 23038 28262 23050 28314
rect 23050 28262 23056 28314
rect 23080 28262 23102 28314
rect 23102 28262 23114 28314
rect 23114 28262 23136 28314
rect 23160 28262 23166 28314
rect 23166 28262 23178 28314
rect 23178 28262 23216 28314
rect 23240 28262 23242 28314
rect 23242 28262 23294 28314
rect 23294 28262 23296 28314
rect 22920 28260 22976 28262
rect 23000 28260 23056 28262
rect 23080 28260 23136 28262
rect 23160 28260 23216 28262
rect 23240 28260 23296 28262
rect 23386 27920 23442 27976
rect 22180 26682 22236 26684
rect 22260 26682 22316 26684
rect 22340 26682 22396 26684
rect 22420 26682 22476 26684
rect 22500 26682 22556 26684
rect 22180 26630 22182 26682
rect 22182 26630 22234 26682
rect 22234 26630 22236 26682
rect 22260 26630 22298 26682
rect 22298 26630 22310 26682
rect 22310 26630 22316 26682
rect 22340 26630 22362 26682
rect 22362 26630 22374 26682
rect 22374 26630 22396 26682
rect 22420 26630 22426 26682
rect 22426 26630 22438 26682
rect 22438 26630 22476 26682
rect 22500 26630 22502 26682
rect 22502 26630 22554 26682
rect 22554 26630 22556 26682
rect 22180 26628 22236 26630
rect 22260 26628 22316 26630
rect 22340 26628 22396 26630
rect 22420 26628 22476 26630
rect 22500 26628 22556 26630
rect 22180 25594 22236 25596
rect 22260 25594 22316 25596
rect 22340 25594 22396 25596
rect 22420 25594 22476 25596
rect 22500 25594 22556 25596
rect 22180 25542 22182 25594
rect 22182 25542 22234 25594
rect 22234 25542 22236 25594
rect 22260 25542 22298 25594
rect 22298 25542 22310 25594
rect 22310 25542 22316 25594
rect 22340 25542 22362 25594
rect 22362 25542 22374 25594
rect 22374 25542 22396 25594
rect 22420 25542 22426 25594
rect 22426 25542 22438 25594
rect 22438 25542 22476 25594
rect 22500 25542 22502 25594
rect 22502 25542 22554 25594
rect 22554 25542 22556 25594
rect 22180 25540 22236 25542
rect 22260 25540 22316 25542
rect 22340 25540 22396 25542
rect 22420 25540 22476 25542
rect 22500 25540 22556 25542
rect 22180 24506 22236 24508
rect 22260 24506 22316 24508
rect 22340 24506 22396 24508
rect 22420 24506 22476 24508
rect 22500 24506 22556 24508
rect 22180 24454 22182 24506
rect 22182 24454 22234 24506
rect 22234 24454 22236 24506
rect 22260 24454 22298 24506
rect 22298 24454 22310 24506
rect 22310 24454 22316 24506
rect 22340 24454 22362 24506
rect 22362 24454 22374 24506
rect 22374 24454 22396 24506
rect 22420 24454 22426 24506
rect 22426 24454 22438 24506
rect 22438 24454 22476 24506
rect 22500 24454 22502 24506
rect 22502 24454 22554 24506
rect 22554 24454 22556 24506
rect 22180 24452 22236 24454
rect 22260 24452 22316 24454
rect 22340 24452 22396 24454
rect 22420 24452 22476 24454
rect 22500 24452 22556 24454
rect 22180 23418 22236 23420
rect 22260 23418 22316 23420
rect 22340 23418 22396 23420
rect 22420 23418 22476 23420
rect 22500 23418 22556 23420
rect 22180 23366 22182 23418
rect 22182 23366 22234 23418
rect 22234 23366 22236 23418
rect 22260 23366 22298 23418
rect 22298 23366 22310 23418
rect 22310 23366 22316 23418
rect 22340 23366 22362 23418
rect 22362 23366 22374 23418
rect 22374 23366 22396 23418
rect 22420 23366 22426 23418
rect 22426 23366 22438 23418
rect 22438 23366 22476 23418
rect 22500 23366 22502 23418
rect 22502 23366 22554 23418
rect 22554 23366 22556 23418
rect 22180 23364 22236 23366
rect 22260 23364 22316 23366
rect 22340 23364 22396 23366
rect 22420 23364 22476 23366
rect 22500 23364 22556 23366
rect 20994 21936 21050 21992
rect 22180 22330 22236 22332
rect 22260 22330 22316 22332
rect 22340 22330 22396 22332
rect 22420 22330 22476 22332
rect 22500 22330 22556 22332
rect 22180 22278 22182 22330
rect 22182 22278 22234 22330
rect 22234 22278 22236 22330
rect 22260 22278 22298 22330
rect 22298 22278 22310 22330
rect 22310 22278 22316 22330
rect 22340 22278 22362 22330
rect 22362 22278 22374 22330
rect 22374 22278 22396 22330
rect 22420 22278 22426 22330
rect 22426 22278 22438 22330
rect 22438 22278 22476 22330
rect 22500 22278 22502 22330
rect 22502 22278 22554 22330
rect 22554 22278 22556 22330
rect 22180 22276 22236 22278
rect 22260 22276 22316 22278
rect 22340 22276 22396 22278
rect 22420 22276 22476 22278
rect 22500 22276 22556 22278
rect 22180 21242 22236 21244
rect 22260 21242 22316 21244
rect 22340 21242 22396 21244
rect 22420 21242 22476 21244
rect 22500 21242 22556 21244
rect 22180 21190 22182 21242
rect 22182 21190 22234 21242
rect 22234 21190 22236 21242
rect 22260 21190 22298 21242
rect 22298 21190 22310 21242
rect 22310 21190 22316 21242
rect 22340 21190 22362 21242
rect 22362 21190 22374 21242
rect 22374 21190 22396 21242
rect 22420 21190 22426 21242
rect 22426 21190 22438 21242
rect 22438 21190 22476 21242
rect 22500 21190 22502 21242
rect 22502 21190 22554 21242
rect 22554 21190 22556 21242
rect 22180 21188 22236 21190
rect 22260 21188 22316 21190
rect 22340 21188 22396 21190
rect 22420 21188 22476 21190
rect 22500 21188 22556 21190
rect 18694 17740 18750 17776
rect 18694 17720 18696 17740
rect 18696 17720 18748 17740
rect 18748 17720 18750 17740
rect 19338 17584 19394 17640
rect 20626 19352 20682 19408
rect 19614 16224 19670 16280
rect 17866 8744 17922 8800
rect 16920 7642 16976 7644
rect 17000 7642 17056 7644
rect 17080 7642 17136 7644
rect 17160 7642 17216 7644
rect 17240 7642 17296 7644
rect 16920 7590 16922 7642
rect 16922 7590 16974 7642
rect 16974 7590 16976 7642
rect 17000 7590 17038 7642
rect 17038 7590 17050 7642
rect 17050 7590 17056 7642
rect 17080 7590 17102 7642
rect 17102 7590 17114 7642
rect 17114 7590 17136 7642
rect 17160 7590 17166 7642
rect 17166 7590 17178 7642
rect 17178 7590 17216 7642
rect 17240 7590 17242 7642
rect 17242 7590 17294 7642
rect 17294 7590 17296 7642
rect 16920 7588 16976 7590
rect 17000 7588 17056 7590
rect 17080 7588 17136 7590
rect 17160 7588 17216 7590
rect 17240 7588 17296 7590
rect 16180 7098 16236 7100
rect 16260 7098 16316 7100
rect 16340 7098 16396 7100
rect 16420 7098 16476 7100
rect 16500 7098 16556 7100
rect 16180 7046 16182 7098
rect 16182 7046 16234 7098
rect 16234 7046 16236 7098
rect 16260 7046 16298 7098
rect 16298 7046 16310 7098
rect 16310 7046 16316 7098
rect 16340 7046 16362 7098
rect 16362 7046 16374 7098
rect 16374 7046 16396 7098
rect 16420 7046 16426 7098
rect 16426 7046 16438 7098
rect 16438 7046 16476 7098
rect 16500 7046 16502 7098
rect 16502 7046 16554 7098
rect 16554 7046 16556 7098
rect 16180 7044 16236 7046
rect 16260 7044 16316 7046
rect 16340 7044 16396 7046
rect 16420 7044 16476 7046
rect 16500 7044 16556 7046
rect 16920 6554 16976 6556
rect 17000 6554 17056 6556
rect 17080 6554 17136 6556
rect 17160 6554 17216 6556
rect 17240 6554 17296 6556
rect 16920 6502 16922 6554
rect 16922 6502 16974 6554
rect 16974 6502 16976 6554
rect 17000 6502 17038 6554
rect 17038 6502 17050 6554
rect 17050 6502 17056 6554
rect 17080 6502 17102 6554
rect 17102 6502 17114 6554
rect 17114 6502 17136 6554
rect 17160 6502 17166 6554
rect 17166 6502 17178 6554
rect 17178 6502 17216 6554
rect 17240 6502 17242 6554
rect 17242 6502 17294 6554
rect 17294 6502 17296 6554
rect 16920 6500 16976 6502
rect 17000 6500 17056 6502
rect 17080 6500 17136 6502
rect 17160 6500 17216 6502
rect 17240 6500 17296 6502
rect 16180 6010 16236 6012
rect 16260 6010 16316 6012
rect 16340 6010 16396 6012
rect 16420 6010 16476 6012
rect 16500 6010 16556 6012
rect 16180 5958 16182 6010
rect 16182 5958 16234 6010
rect 16234 5958 16236 6010
rect 16260 5958 16298 6010
rect 16298 5958 16310 6010
rect 16310 5958 16316 6010
rect 16340 5958 16362 6010
rect 16362 5958 16374 6010
rect 16374 5958 16396 6010
rect 16420 5958 16426 6010
rect 16426 5958 16438 6010
rect 16438 5958 16476 6010
rect 16500 5958 16502 6010
rect 16502 5958 16554 6010
rect 16554 5958 16556 6010
rect 16180 5956 16236 5958
rect 16260 5956 16316 5958
rect 16340 5956 16396 5958
rect 16420 5956 16476 5958
rect 16500 5956 16556 5958
rect 16920 5466 16976 5468
rect 17000 5466 17056 5468
rect 17080 5466 17136 5468
rect 17160 5466 17216 5468
rect 17240 5466 17296 5468
rect 16920 5414 16922 5466
rect 16922 5414 16974 5466
rect 16974 5414 16976 5466
rect 17000 5414 17038 5466
rect 17038 5414 17050 5466
rect 17050 5414 17056 5466
rect 17080 5414 17102 5466
rect 17102 5414 17114 5466
rect 17114 5414 17136 5466
rect 17160 5414 17166 5466
rect 17166 5414 17178 5466
rect 17178 5414 17216 5466
rect 17240 5414 17242 5466
rect 17242 5414 17294 5466
rect 17294 5414 17296 5466
rect 16920 5412 16976 5414
rect 17000 5412 17056 5414
rect 17080 5412 17136 5414
rect 17160 5412 17216 5414
rect 17240 5412 17296 5414
rect 16180 4922 16236 4924
rect 16260 4922 16316 4924
rect 16340 4922 16396 4924
rect 16420 4922 16476 4924
rect 16500 4922 16556 4924
rect 16180 4870 16182 4922
rect 16182 4870 16234 4922
rect 16234 4870 16236 4922
rect 16260 4870 16298 4922
rect 16298 4870 16310 4922
rect 16310 4870 16316 4922
rect 16340 4870 16362 4922
rect 16362 4870 16374 4922
rect 16374 4870 16396 4922
rect 16420 4870 16426 4922
rect 16426 4870 16438 4922
rect 16438 4870 16476 4922
rect 16500 4870 16502 4922
rect 16502 4870 16554 4922
rect 16554 4870 16556 4922
rect 16180 4868 16236 4870
rect 16260 4868 16316 4870
rect 16340 4868 16396 4870
rect 16420 4868 16476 4870
rect 16500 4868 16556 4870
rect 16920 4378 16976 4380
rect 17000 4378 17056 4380
rect 17080 4378 17136 4380
rect 17160 4378 17216 4380
rect 17240 4378 17296 4380
rect 16920 4326 16922 4378
rect 16922 4326 16974 4378
rect 16974 4326 16976 4378
rect 17000 4326 17038 4378
rect 17038 4326 17050 4378
rect 17050 4326 17056 4378
rect 17080 4326 17102 4378
rect 17102 4326 17114 4378
rect 17114 4326 17136 4378
rect 17160 4326 17166 4378
rect 17166 4326 17178 4378
rect 17178 4326 17216 4378
rect 17240 4326 17242 4378
rect 17242 4326 17294 4378
rect 17294 4326 17296 4378
rect 16920 4324 16976 4326
rect 17000 4324 17056 4326
rect 17080 4324 17136 4326
rect 17160 4324 17216 4326
rect 17240 4324 17296 4326
rect 16180 3834 16236 3836
rect 16260 3834 16316 3836
rect 16340 3834 16396 3836
rect 16420 3834 16476 3836
rect 16500 3834 16556 3836
rect 16180 3782 16182 3834
rect 16182 3782 16234 3834
rect 16234 3782 16236 3834
rect 16260 3782 16298 3834
rect 16298 3782 16310 3834
rect 16310 3782 16316 3834
rect 16340 3782 16362 3834
rect 16362 3782 16374 3834
rect 16374 3782 16396 3834
rect 16420 3782 16426 3834
rect 16426 3782 16438 3834
rect 16438 3782 16476 3834
rect 16500 3782 16502 3834
rect 16502 3782 16554 3834
rect 16554 3782 16556 3834
rect 16180 3780 16236 3782
rect 16260 3780 16316 3782
rect 16340 3780 16396 3782
rect 16420 3780 16476 3782
rect 16500 3780 16556 3782
rect 16920 3290 16976 3292
rect 17000 3290 17056 3292
rect 17080 3290 17136 3292
rect 17160 3290 17216 3292
rect 17240 3290 17296 3292
rect 16920 3238 16922 3290
rect 16922 3238 16974 3290
rect 16974 3238 16976 3290
rect 17000 3238 17038 3290
rect 17038 3238 17050 3290
rect 17050 3238 17056 3290
rect 17080 3238 17102 3290
rect 17102 3238 17114 3290
rect 17114 3238 17136 3290
rect 17160 3238 17166 3290
rect 17166 3238 17178 3290
rect 17178 3238 17216 3290
rect 17240 3238 17242 3290
rect 17242 3238 17294 3290
rect 17294 3238 17296 3290
rect 16920 3236 16976 3238
rect 17000 3236 17056 3238
rect 17080 3236 17136 3238
rect 17160 3236 17216 3238
rect 17240 3236 17296 3238
rect 22180 20154 22236 20156
rect 22260 20154 22316 20156
rect 22340 20154 22396 20156
rect 22420 20154 22476 20156
rect 22500 20154 22556 20156
rect 22180 20102 22182 20154
rect 22182 20102 22234 20154
rect 22234 20102 22236 20154
rect 22260 20102 22298 20154
rect 22298 20102 22310 20154
rect 22310 20102 22316 20154
rect 22340 20102 22362 20154
rect 22362 20102 22374 20154
rect 22374 20102 22396 20154
rect 22420 20102 22426 20154
rect 22426 20102 22438 20154
rect 22438 20102 22476 20154
rect 22500 20102 22502 20154
rect 22502 20102 22554 20154
rect 22554 20102 22556 20154
rect 22180 20100 22236 20102
rect 22260 20100 22316 20102
rect 22340 20100 22396 20102
rect 22420 20100 22476 20102
rect 22500 20100 22556 20102
rect 21086 17584 21142 17640
rect 20994 16224 21050 16280
rect 22180 19066 22236 19068
rect 22260 19066 22316 19068
rect 22340 19066 22396 19068
rect 22420 19066 22476 19068
rect 22500 19066 22556 19068
rect 22180 19014 22182 19066
rect 22182 19014 22234 19066
rect 22234 19014 22236 19066
rect 22260 19014 22298 19066
rect 22298 19014 22310 19066
rect 22310 19014 22316 19066
rect 22340 19014 22362 19066
rect 22362 19014 22374 19066
rect 22374 19014 22396 19066
rect 22420 19014 22426 19066
rect 22426 19014 22438 19066
rect 22438 19014 22476 19066
rect 22500 19014 22502 19066
rect 22502 19014 22554 19066
rect 22554 19014 22556 19066
rect 22180 19012 22236 19014
rect 22260 19012 22316 19014
rect 22340 19012 22396 19014
rect 22420 19012 22476 19014
rect 22500 19012 22556 19014
rect 22180 17978 22236 17980
rect 22260 17978 22316 17980
rect 22340 17978 22396 17980
rect 22420 17978 22476 17980
rect 22500 17978 22556 17980
rect 22180 17926 22182 17978
rect 22182 17926 22234 17978
rect 22234 17926 22236 17978
rect 22260 17926 22298 17978
rect 22298 17926 22310 17978
rect 22310 17926 22316 17978
rect 22340 17926 22362 17978
rect 22362 17926 22374 17978
rect 22374 17926 22396 17978
rect 22420 17926 22426 17978
rect 22426 17926 22438 17978
rect 22438 17926 22476 17978
rect 22500 17926 22502 17978
rect 22502 17926 22554 17978
rect 22554 17926 22556 17978
rect 22180 17924 22236 17926
rect 22260 17924 22316 17926
rect 22340 17924 22396 17926
rect 22420 17924 22476 17926
rect 22500 17924 22556 17926
rect 22180 16890 22236 16892
rect 22260 16890 22316 16892
rect 22340 16890 22396 16892
rect 22420 16890 22476 16892
rect 22500 16890 22556 16892
rect 22180 16838 22182 16890
rect 22182 16838 22234 16890
rect 22234 16838 22236 16890
rect 22260 16838 22298 16890
rect 22298 16838 22310 16890
rect 22310 16838 22316 16890
rect 22340 16838 22362 16890
rect 22362 16838 22374 16890
rect 22374 16838 22396 16890
rect 22420 16838 22426 16890
rect 22426 16838 22438 16890
rect 22438 16838 22476 16890
rect 22500 16838 22502 16890
rect 22502 16838 22554 16890
rect 22554 16838 22556 16890
rect 22180 16836 22236 16838
rect 22260 16836 22316 16838
rect 22340 16836 22396 16838
rect 22420 16836 22476 16838
rect 22500 16836 22556 16838
rect 22180 15802 22236 15804
rect 22260 15802 22316 15804
rect 22340 15802 22396 15804
rect 22420 15802 22476 15804
rect 22500 15802 22556 15804
rect 22180 15750 22182 15802
rect 22182 15750 22234 15802
rect 22234 15750 22236 15802
rect 22260 15750 22298 15802
rect 22298 15750 22310 15802
rect 22310 15750 22316 15802
rect 22340 15750 22362 15802
rect 22362 15750 22374 15802
rect 22374 15750 22396 15802
rect 22420 15750 22426 15802
rect 22426 15750 22438 15802
rect 22438 15750 22476 15802
rect 22500 15750 22502 15802
rect 22502 15750 22554 15802
rect 22554 15750 22556 15802
rect 22180 15748 22236 15750
rect 22260 15748 22316 15750
rect 22340 15748 22396 15750
rect 22420 15748 22476 15750
rect 22500 15748 22556 15750
rect 22180 14714 22236 14716
rect 22260 14714 22316 14716
rect 22340 14714 22396 14716
rect 22420 14714 22476 14716
rect 22500 14714 22556 14716
rect 22180 14662 22182 14714
rect 22182 14662 22234 14714
rect 22234 14662 22236 14714
rect 22260 14662 22298 14714
rect 22298 14662 22310 14714
rect 22310 14662 22316 14714
rect 22340 14662 22362 14714
rect 22362 14662 22374 14714
rect 22374 14662 22396 14714
rect 22420 14662 22426 14714
rect 22426 14662 22438 14714
rect 22438 14662 22476 14714
rect 22500 14662 22502 14714
rect 22502 14662 22554 14714
rect 22554 14662 22556 14714
rect 22180 14660 22236 14662
rect 22260 14660 22316 14662
rect 22340 14660 22396 14662
rect 22420 14660 22476 14662
rect 22500 14660 22556 14662
rect 22920 27226 22976 27228
rect 23000 27226 23056 27228
rect 23080 27226 23136 27228
rect 23160 27226 23216 27228
rect 23240 27226 23296 27228
rect 22920 27174 22922 27226
rect 22922 27174 22974 27226
rect 22974 27174 22976 27226
rect 23000 27174 23038 27226
rect 23038 27174 23050 27226
rect 23050 27174 23056 27226
rect 23080 27174 23102 27226
rect 23102 27174 23114 27226
rect 23114 27174 23136 27226
rect 23160 27174 23166 27226
rect 23166 27174 23178 27226
rect 23178 27174 23216 27226
rect 23240 27174 23242 27226
rect 23242 27174 23294 27226
rect 23294 27174 23296 27226
rect 22920 27172 22976 27174
rect 23000 27172 23056 27174
rect 23080 27172 23136 27174
rect 23160 27172 23216 27174
rect 23240 27172 23296 27174
rect 22920 26138 22976 26140
rect 23000 26138 23056 26140
rect 23080 26138 23136 26140
rect 23160 26138 23216 26140
rect 23240 26138 23296 26140
rect 22920 26086 22922 26138
rect 22922 26086 22974 26138
rect 22974 26086 22976 26138
rect 23000 26086 23038 26138
rect 23038 26086 23050 26138
rect 23050 26086 23056 26138
rect 23080 26086 23102 26138
rect 23102 26086 23114 26138
rect 23114 26086 23136 26138
rect 23160 26086 23166 26138
rect 23166 26086 23178 26138
rect 23178 26086 23216 26138
rect 23240 26086 23242 26138
rect 23242 26086 23294 26138
rect 23294 26086 23296 26138
rect 22920 26084 22976 26086
rect 23000 26084 23056 26086
rect 23080 26084 23136 26086
rect 23160 26084 23216 26086
rect 23240 26084 23296 26086
rect 22920 25050 22976 25052
rect 23000 25050 23056 25052
rect 23080 25050 23136 25052
rect 23160 25050 23216 25052
rect 23240 25050 23296 25052
rect 22920 24998 22922 25050
rect 22922 24998 22974 25050
rect 22974 24998 22976 25050
rect 23000 24998 23038 25050
rect 23038 24998 23050 25050
rect 23050 24998 23056 25050
rect 23080 24998 23102 25050
rect 23102 24998 23114 25050
rect 23114 24998 23136 25050
rect 23160 24998 23166 25050
rect 23166 24998 23178 25050
rect 23178 24998 23216 25050
rect 23240 24998 23242 25050
rect 23242 24998 23294 25050
rect 23294 24998 23296 25050
rect 22920 24996 22976 24998
rect 23000 24996 23056 24998
rect 23080 24996 23136 24998
rect 23160 24996 23216 24998
rect 23240 24996 23296 24998
rect 22920 23962 22976 23964
rect 23000 23962 23056 23964
rect 23080 23962 23136 23964
rect 23160 23962 23216 23964
rect 23240 23962 23296 23964
rect 22920 23910 22922 23962
rect 22922 23910 22974 23962
rect 22974 23910 22976 23962
rect 23000 23910 23038 23962
rect 23038 23910 23050 23962
rect 23050 23910 23056 23962
rect 23080 23910 23102 23962
rect 23102 23910 23114 23962
rect 23114 23910 23136 23962
rect 23160 23910 23166 23962
rect 23166 23910 23178 23962
rect 23178 23910 23216 23962
rect 23240 23910 23242 23962
rect 23242 23910 23294 23962
rect 23294 23910 23296 23962
rect 22920 23908 22976 23910
rect 23000 23908 23056 23910
rect 23080 23908 23136 23910
rect 23160 23908 23216 23910
rect 23240 23908 23296 23910
rect 22920 22874 22976 22876
rect 23000 22874 23056 22876
rect 23080 22874 23136 22876
rect 23160 22874 23216 22876
rect 23240 22874 23296 22876
rect 22920 22822 22922 22874
rect 22922 22822 22974 22874
rect 22974 22822 22976 22874
rect 23000 22822 23038 22874
rect 23038 22822 23050 22874
rect 23050 22822 23056 22874
rect 23080 22822 23102 22874
rect 23102 22822 23114 22874
rect 23114 22822 23136 22874
rect 23160 22822 23166 22874
rect 23166 22822 23178 22874
rect 23178 22822 23216 22874
rect 23240 22822 23242 22874
rect 23242 22822 23294 22874
rect 23294 22822 23296 22874
rect 22920 22820 22976 22822
rect 23000 22820 23056 22822
rect 23080 22820 23136 22822
rect 23160 22820 23216 22822
rect 23240 22820 23296 22822
rect 22920 21786 22976 21788
rect 23000 21786 23056 21788
rect 23080 21786 23136 21788
rect 23160 21786 23216 21788
rect 23240 21786 23296 21788
rect 22920 21734 22922 21786
rect 22922 21734 22974 21786
rect 22974 21734 22976 21786
rect 23000 21734 23038 21786
rect 23038 21734 23050 21786
rect 23050 21734 23056 21786
rect 23080 21734 23102 21786
rect 23102 21734 23114 21786
rect 23114 21734 23136 21786
rect 23160 21734 23166 21786
rect 23166 21734 23178 21786
rect 23178 21734 23216 21786
rect 23240 21734 23242 21786
rect 23242 21734 23294 21786
rect 23294 21734 23296 21786
rect 22920 21732 22976 21734
rect 23000 21732 23056 21734
rect 23080 21732 23136 21734
rect 23160 21732 23216 21734
rect 23240 21732 23296 21734
rect 22920 20698 22976 20700
rect 23000 20698 23056 20700
rect 23080 20698 23136 20700
rect 23160 20698 23216 20700
rect 23240 20698 23296 20700
rect 22920 20646 22922 20698
rect 22922 20646 22974 20698
rect 22974 20646 22976 20698
rect 23000 20646 23038 20698
rect 23038 20646 23050 20698
rect 23050 20646 23056 20698
rect 23080 20646 23102 20698
rect 23102 20646 23114 20698
rect 23114 20646 23136 20698
rect 23160 20646 23166 20698
rect 23166 20646 23178 20698
rect 23178 20646 23216 20698
rect 23240 20646 23242 20698
rect 23242 20646 23294 20698
rect 23294 20646 23296 20698
rect 22920 20644 22976 20646
rect 23000 20644 23056 20646
rect 23080 20644 23136 20646
rect 23160 20644 23216 20646
rect 23240 20644 23296 20646
rect 22920 19610 22976 19612
rect 23000 19610 23056 19612
rect 23080 19610 23136 19612
rect 23160 19610 23216 19612
rect 23240 19610 23296 19612
rect 22920 19558 22922 19610
rect 22922 19558 22974 19610
rect 22974 19558 22976 19610
rect 23000 19558 23038 19610
rect 23038 19558 23050 19610
rect 23050 19558 23056 19610
rect 23080 19558 23102 19610
rect 23102 19558 23114 19610
rect 23114 19558 23136 19610
rect 23160 19558 23166 19610
rect 23166 19558 23178 19610
rect 23178 19558 23216 19610
rect 23240 19558 23242 19610
rect 23242 19558 23294 19610
rect 23294 19558 23296 19610
rect 22920 19556 22976 19558
rect 23000 19556 23056 19558
rect 23080 19556 23136 19558
rect 23160 19556 23216 19558
rect 23240 19556 23296 19558
rect 22920 18522 22976 18524
rect 23000 18522 23056 18524
rect 23080 18522 23136 18524
rect 23160 18522 23216 18524
rect 23240 18522 23296 18524
rect 22920 18470 22922 18522
rect 22922 18470 22974 18522
rect 22974 18470 22976 18522
rect 23000 18470 23038 18522
rect 23038 18470 23050 18522
rect 23050 18470 23056 18522
rect 23080 18470 23102 18522
rect 23102 18470 23114 18522
rect 23114 18470 23136 18522
rect 23160 18470 23166 18522
rect 23166 18470 23178 18522
rect 23178 18470 23216 18522
rect 23240 18470 23242 18522
rect 23242 18470 23294 18522
rect 23294 18470 23296 18522
rect 22920 18468 22976 18470
rect 23000 18468 23056 18470
rect 23080 18468 23136 18470
rect 23160 18468 23216 18470
rect 23240 18468 23296 18470
rect 22920 17434 22976 17436
rect 23000 17434 23056 17436
rect 23080 17434 23136 17436
rect 23160 17434 23216 17436
rect 23240 17434 23296 17436
rect 22920 17382 22922 17434
rect 22922 17382 22974 17434
rect 22974 17382 22976 17434
rect 23000 17382 23038 17434
rect 23038 17382 23050 17434
rect 23050 17382 23056 17434
rect 23080 17382 23102 17434
rect 23102 17382 23114 17434
rect 23114 17382 23136 17434
rect 23160 17382 23166 17434
rect 23166 17382 23178 17434
rect 23178 17382 23216 17434
rect 23240 17382 23242 17434
rect 23242 17382 23294 17434
rect 23294 17382 23296 17434
rect 22920 17380 22976 17382
rect 23000 17380 23056 17382
rect 23080 17380 23136 17382
rect 23160 17380 23216 17382
rect 23240 17380 23296 17382
rect 22920 16346 22976 16348
rect 23000 16346 23056 16348
rect 23080 16346 23136 16348
rect 23160 16346 23216 16348
rect 23240 16346 23296 16348
rect 22920 16294 22922 16346
rect 22922 16294 22974 16346
rect 22974 16294 22976 16346
rect 23000 16294 23038 16346
rect 23038 16294 23050 16346
rect 23050 16294 23056 16346
rect 23080 16294 23102 16346
rect 23102 16294 23114 16346
rect 23114 16294 23136 16346
rect 23160 16294 23166 16346
rect 23166 16294 23178 16346
rect 23178 16294 23216 16346
rect 23240 16294 23242 16346
rect 23242 16294 23294 16346
rect 23294 16294 23296 16346
rect 22920 16292 22976 16294
rect 23000 16292 23056 16294
rect 23080 16292 23136 16294
rect 23160 16292 23216 16294
rect 23240 16292 23296 16294
rect 22920 15258 22976 15260
rect 23000 15258 23056 15260
rect 23080 15258 23136 15260
rect 23160 15258 23216 15260
rect 23240 15258 23296 15260
rect 22920 15206 22922 15258
rect 22922 15206 22974 15258
rect 22974 15206 22976 15258
rect 23000 15206 23038 15258
rect 23038 15206 23050 15258
rect 23050 15206 23056 15258
rect 23080 15206 23102 15258
rect 23102 15206 23114 15258
rect 23114 15206 23136 15258
rect 23160 15206 23166 15258
rect 23166 15206 23178 15258
rect 23178 15206 23216 15258
rect 23240 15206 23242 15258
rect 23242 15206 23294 15258
rect 23294 15206 23296 15258
rect 22920 15204 22976 15206
rect 23000 15204 23056 15206
rect 23080 15204 23136 15206
rect 23160 15204 23216 15206
rect 23240 15204 23296 15206
rect 22180 13626 22236 13628
rect 22260 13626 22316 13628
rect 22340 13626 22396 13628
rect 22420 13626 22476 13628
rect 22500 13626 22556 13628
rect 22180 13574 22182 13626
rect 22182 13574 22234 13626
rect 22234 13574 22236 13626
rect 22260 13574 22298 13626
rect 22298 13574 22310 13626
rect 22310 13574 22316 13626
rect 22340 13574 22362 13626
rect 22362 13574 22374 13626
rect 22374 13574 22396 13626
rect 22420 13574 22426 13626
rect 22426 13574 22438 13626
rect 22438 13574 22476 13626
rect 22500 13574 22502 13626
rect 22502 13574 22554 13626
rect 22554 13574 22556 13626
rect 22180 13572 22236 13574
rect 22260 13572 22316 13574
rect 22340 13572 22396 13574
rect 22420 13572 22476 13574
rect 22500 13572 22556 13574
rect 22180 12538 22236 12540
rect 22260 12538 22316 12540
rect 22340 12538 22396 12540
rect 22420 12538 22476 12540
rect 22500 12538 22556 12540
rect 22180 12486 22182 12538
rect 22182 12486 22234 12538
rect 22234 12486 22236 12538
rect 22260 12486 22298 12538
rect 22298 12486 22310 12538
rect 22310 12486 22316 12538
rect 22340 12486 22362 12538
rect 22362 12486 22374 12538
rect 22374 12486 22396 12538
rect 22420 12486 22426 12538
rect 22426 12486 22438 12538
rect 22438 12486 22476 12538
rect 22500 12486 22502 12538
rect 22502 12486 22554 12538
rect 22554 12486 22556 12538
rect 22180 12484 22236 12486
rect 22260 12484 22316 12486
rect 22340 12484 22396 12486
rect 22420 12484 22476 12486
rect 22500 12484 22556 12486
rect 22180 11450 22236 11452
rect 22260 11450 22316 11452
rect 22340 11450 22396 11452
rect 22420 11450 22476 11452
rect 22500 11450 22556 11452
rect 22180 11398 22182 11450
rect 22182 11398 22234 11450
rect 22234 11398 22236 11450
rect 22260 11398 22298 11450
rect 22298 11398 22310 11450
rect 22310 11398 22316 11450
rect 22340 11398 22362 11450
rect 22362 11398 22374 11450
rect 22374 11398 22396 11450
rect 22420 11398 22426 11450
rect 22426 11398 22438 11450
rect 22438 11398 22476 11450
rect 22500 11398 22502 11450
rect 22502 11398 22554 11450
rect 22554 11398 22556 11450
rect 22180 11396 22236 11398
rect 22260 11396 22316 11398
rect 22340 11396 22396 11398
rect 22420 11396 22476 11398
rect 22500 11396 22556 11398
rect 22180 10362 22236 10364
rect 22260 10362 22316 10364
rect 22340 10362 22396 10364
rect 22420 10362 22476 10364
rect 22500 10362 22556 10364
rect 22180 10310 22182 10362
rect 22182 10310 22234 10362
rect 22234 10310 22236 10362
rect 22260 10310 22298 10362
rect 22298 10310 22310 10362
rect 22310 10310 22316 10362
rect 22340 10310 22362 10362
rect 22362 10310 22374 10362
rect 22374 10310 22396 10362
rect 22420 10310 22426 10362
rect 22426 10310 22438 10362
rect 22438 10310 22476 10362
rect 22500 10310 22502 10362
rect 22502 10310 22554 10362
rect 22554 10310 22556 10362
rect 22180 10308 22236 10310
rect 22260 10308 22316 10310
rect 22340 10308 22396 10310
rect 22420 10308 22476 10310
rect 22500 10308 22556 10310
rect 22558 9696 22614 9752
rect 22920 14170 22976 14172
rect 23000 14170 23056 14172
rect 23080 14170 23136 14172
rect 23160 14170 23216 14172
rect 23240 14170 23296 14172
rect 22920 14118 22922 14170
rect 22922 14118 22974 14170
rect 22974 14118 22976 14170
rect 23000 14118 23038 14170
rect 23038 14118 23050 14170
rect 23050 14118 23056 14170
rect 23080 14118 23102 14170
rect 23102 14118 23114 14170
rect 23114 14118 23136 14170
rect 23160 14118 23166 14170
rect 23166 14118 23178 14170
rect 23178 14118 23216 14170
rect 23240 14118 23242 14170
rect 23242 14118 23294 14170
rect 23294 14118 23296 14170
rect 22920 14116 22976 14118
rect 23000 14116 23056 14118
rect 23080 14116 23136 14118
rect 23160 14116 23216 14118
rect 23240 14116 23296 14118
rect 22920 13082 22976 13084
rect 23000 13082 23056 13084
rect 23080 13082 23136 13084
rect 23160 13082 23216 13084
rect 23240 13082 23296 13084
rect 22920 13030 22922 13082
rect 22922 13030 22974 13082
rect 22974 13030 22976 13082
rect 23000 13030 23038 13082
rect 23038 13030 23050 13082
rect 23050 13030 23056 13082
rect 23080 13030 23102 13082
rect 23102 13030 23114 13082
rect 23114 13030 23136 13082
rect 23160 13030 23166 13082
rect 23166 13030 23178 13082
rect 23178 13030 23216 13082
rect 23240 13030 23242 13082
rect 23242 13030 23294 13082
rect 23294 13030 23296 13082
rect 22920 13028 22976 13030
rect 23000 13028 23056 13030
rect 23080 13028 23136 13030
rect 23160 13028 23216 13030
rect 23240 13028 23296 13030
rect 28920 31578 28976 31580
rect 29000 31578 29056 31580
rect 29080 31578 29136 31580
rect 29160 31578 29216 31580
rect 29240 31578 29296 31580
rect 28920 31526 28922 31578
rect 28922 31526 28974 31578
rect 28974 31526 28976 31578
rect 29000 31526 29038 31578
rect 29038 31526 29050 31578
rect 29050 31526 29056 31578
rect 29080 31526 29102 31578
rect 29102 31526 29114 31578
rect 29114 31526 29136 31578
rect 29160 31526 29166 31578
rect 29166 31526 29178 31578
rect 29178 31526 29216 31578
rect 29240 31526 29242 31578
rect 29242 31526 29294 31578
rect 29294 31526 29296 31578
rect 28920 31524 28976 31526
rect 29000 31524 29056 31526
rect 29080 31524 29136 31526
rect 29160 31524 29216 31526
rect 29240 31524 29296 31526
rect 28180 31034 28236 31036
rect 28260 31034 28316 31036
rect 28340 31034 28396 31036
rect 28420 31034 28476 31036
rect 28500 31034 28556 31036
rect 28180 30982 28182 31034
rect 28182 30982 28234 31034
rect 28234 30982 28236 31034
rect 28260 30982 28298 31034
rect 28298 30982 28310 31034
rect 28310 30982 28316 31034
rect 28340 30982 28362 31034
rect 28362 30982 28374 31034
rect 28374 30982 28396 31034
rect 28420 30982 28426 31034
rect 28426 30982 28438 31034
rect 28438 30982 28476 31034
rect 28500 30982 28502 31034
rect 28502 30982 28554 31034
rect 28554 30982 28556 31034
rect 28180 30980 28236 30982
rect 28260 30980 28316 30982
rect 28340 30980 28396 30982
rect 28420 30980 28476 30982
rect 28500 30980 28556 30982
rect 24030 27648 24086 27704
rect 24490 19932 24492 19952
rect 24492 19932 24544 19952
rect 24544 19932 24546 19952
rect 24490 19896 24546 19932
rect 23202 12144 23258 12200
rect 22920 11994 22976 11996
rect 23000 11994 23056 11996
rect 23080 11994 23136 11996
rect 23160 11994 23216 11996
rect 23240 11994 23296 11996
rect 22920 11942 22922 11994
rect 22922 11942 22974 11994
rect 22974 11942 22976 11994
rect 23000 11942 23038 11994
rect 23038 11942 23050 11994
rect 23050 11942 23056 11994
rect 23080 11942 23102 11994
rect 23102 11942 23114 11994
rect 23114 11942 23136 11994
rect 23160 11942 23166 11994
rect 23166 11942 23178 11994
rect 23178 11942 23216 11994
rect 23240 11942 23242 11994
rect 23242 11942 23294 11994
rect 23294 11942 23296 11994
rect 22920 11940 22976 11942
rect 23000 11940 23056 11942
rect 23080 11940 23136 11942
rect 23160 11940 23216 11942
rect 23240 11940 23296 11942
rect 23570 11872 23626 11928
rect 22920 10906 22976 10908
rect 23000 10906 23056 10908
rect 23080 10906 23136 10908
rect 23160 10906 23216 10908
rect 23240 10906 23296 10908
rect 22920 10854 22922 10906
rect 22922 10854 22974 10906
rect 22974 10854 22976 10906
rect 23000 10854 23038 10906
rect 23038 10854 23050 10906
rect 23050 10854 23056 10906
rect 23080 10854 23102 10906
rect 23102 10854 23114 10906
rect 23114 10854 23136 10906
rect 23160 10854 23166 10906
rect 23166 10854 23178 10906
rect 23178 10854 23216 10906
rect 23240 10854 23242 10906
rect 23242 10854 23294 10906
rect 23294 10854 23296 10906
rect 22920 10852 22976 10854
rect 23000 10852 23056 10854
rect 23080 10852 23136 10854
rect 23160 10852 23216 10854
rect 23240 10852 23296 10854
rect 23018 9968 23074 10024
rect 22742 9632 22798 9688
rect 22180 9274 22236 9276
rect 22260 9274 22316 9276
rect 22340 9274 22396 9276
rect 22420 9274 22476 9276
rect 22500 9274 22556 9276
rect 22180 9222 22182 9274
rect 22182 9222 22234 9274
rect 22234 9222 22236 9274
rect 22260 9222 22298 9274
rect 22298 9222 22310 9274
rect 22310 9222 22316 9274
rect 22340 9222 22362 9274
rect 22362 9222 22374 9274
rect 22374 9222 22396 9274
rect 22420 9222 22426 9274
rect 22426 9222 22438 9274
rect 22438 9222 22476 9274
rect 22500 9222 22502 9274
rect 22502 9222 22554 9274
rect 22554 9222 22556 9274
rect 22180 9220 22236 9222
rect 22260 9220 22316 9222
rect 22340 9220 22396 9222
rect 22420 9220 22476 9222
rect 22500 9220 22556 9222
rect 22180 8186 22236 8188
rect 22260 8186 22316 8188
rect 22340 8186 22396 8188
rect 22420 8186 22476 8188
rect 22500 8186 22556 8188
rect 22180 8134 22182 8186
rect 22182 8134 22234 8186
rect 22234 8134 22236 8186
rect 22260 8134 22298 8186
rect 22298 8134 22310 8186
rect 22310 8134 22316 8186
rect 22340 8134 22362 8186
rect 22362 8134 22374 8186
rect 22374 8134 22396 8186
rect 22420 8134 22426 8186
rect 22426 8134 22438 8186
rect 22438 8134 22476 8186
rect 22500 8134 22502 8186
rect 22502 8134 22554 8186
rect 22554 8134 22556 8186
rect 22180 8132 22236 8134
rect 22260 8132 22316 8134
rect 22340 8132 22396 8134
rect 22420 8132 22476 8134
rect 22500 8132 22556 8134
rect 22180 7098 22236 7100
rect 22260 7098 22316 7100
rect 22340 7098 22396 7100
rect 22420 7098 22476 7100
rect 22500 7098 22556 7100
rect 22180 7046 22182 7098
rect 22182 7046 22234 7098
rect 22234 7046 22236 7098
rect 22260 7046 22298 7098
rect 22298 7046 22310 7098
rect 22310 7046 22316 7098
rect 22340 7046 22362 7098
rect 22362 7046 22374 7098
rect 22374 7046 22396 7098
rect 22420 7046 22426 7098
rect 22426 7046 22438 7098
rect 22438 7046 22476 7098
rect 22500 7046 22502 7098
rect 22502 7046 22554 7098
rect 22554 7046 22556 7098
rect 22180 7044 22236 7046
rect 22260 7044 22316 7046
rect 22340 7044 22396 7046
rect 22420 7044 22476 7046
rect 22500 7044 22556 7046
rect 22920 9818 22976 9820
rect 23000 9818 23056 9820
rect 23080 9818 23136 9820
rect 23160 9818 23216 9820
rect 23240 9818 23296 9820
rect 22920 9766 22922 9818
rect 22922 9766 22974 9818
rect 22974 9766 22976 9818
rect 23000 9766 23038 9818
rect 23038 9766 23050 9818
rect 23050 9766 23056 9818
rect 23080 9766 23102 9818
rect 23102 9766 23114 9818
rect 23114 9766 23136 9818
rect 23160 9766 23166 9818
rect 23166 9766 23178 9818
rect 23178 9766 23216 9818
rect 23240 9766 23242 9818
rect 23242 9766 23294 9818
rect 23294 9766 23296 9818
rect 22920 9764 22976 9766
rect 23000 9764 23056 9766
rect 23080 9764 23136 9766
rect 23160 9764 23216 9766
rect 23240 9764 23296 9766
rect 23294 9632 23350 9688
rect 23294 8880 23350 8936
rect 22920 8730 22976 8732
rect 23000 8730 23056 8732
rect 23080 8730 23136 8732
rect 23160 8730 23216 8732
rect 23240 8730 23296 8732
rect 22920 8678 22922 8730
rect 22922 8678 22974 8730
rect 22974 8678 22976 8730
rect 23000 8678 23038 8730
rect 23038 8678 23050 8730
rect 23050 8678 23056 8730
rect 23080 8678 23102 8730
rect 23102 8678 23114 8730
rect 23114 8678 23136 8730
rect 23160 8678 23166 8730
rect 23166 8678 23178 8730
rect 23178 8678 23216 8730
rect 23240 8678 23242 8730
rect 23242 8678 23294 8730
rect 23294 8678 23296 8730
rect 22920 8676 22976 8678
rect 23000 8676 23056 8678
rect 23080 8676 23136 8678
rect 23160 8676 23216 8678
rect 23240 8676 23296 8678
rect 22920 7642 22976 7644
rect 23000 7642 23056 7644
rect 23080 7642 23136 7644
rect 23160 7642 23216 7644
rect 23240 7642 23296 7644
rect 22920 7590 22922 7642
rect 22922 7590 22974 7642
rect 22974 7590 22976 7642
rect 23000 7590 23038 7642
rect 23038 7590 23050 7642
rect 23050 7590 23056 7642
rect 23080 7590 23102 7642
rect 23102 7590 23114 7642
rect 23114 7590 23136 7642
rect 23160 7590 23166 7642
rect 23166 7590 23178 7642
rect 23178 7590 23216 7642
rect 23240 7590 23242 7642
rect 23242 7590 23294 7642
rect 23294 7590 23296 7642
rect 22920 7588 22976 7590
rect 23000 7588 23056 7590
rect 23080 7588 23136 7590
rect 23160 7588 23216 7590
rect 23240 7588 23296 7590
rect 22920 6554 22976 6556
rect 23000 6554 23056 6556
rect 23080 6554 23136 6556
rect 23160 6554 23216 6556
rect 23240 6554 23296 6556
rect 22920 6502 22922 6554
rect 22922 6502 22974 6554
rect 22974 6502 22976 6554
rect 23000 6502 23038 6554
rect 23038 6502 23050 6554
rect 23050 6502 23056 6554
rect 23080 6502 23102 6554
rect 23102 6502 23114 6554
rect 23114 6502 23136 6554
rect 23160 6502 23166 6554
rect 23166 6502 23178 6554
rect 23178 6502 23216 6554
rect 23240 6502 23242 6554
rect 23242 6502 23294 6554
rect 23294 6502 23296 6554
rect 22920 6500 22976 6502
rect 23000 6500 23056 6502
rect 23080 6500 23136 6502
rect 23160 6500 23216 6502
rect 23240 6500 23296 6502
rect 22180 6010 22236 6012
rect 22260 6010 22316 6012
rect 22340 6010 22396 6012
rect 22420 6010 22476 6012
rect 22500 6010 22556 6012
rect 22180 5958 22182 6010
rect 22182 5958 22234 6010
rect 22234 5958 22236 6010
rect 22260 5958 22298 6010
rect 22298 5958 22310 6010
rect 22310 5958 22316 6010
rect 22340 5958 22362 6010
rect 22362 5958 22374 6010
rect 22374 5958 22396 6010
rect 22420 5958 22426 6010
rect 22426 5958 22438 6010
rect 22438 5958 22476 6010
rect 22500 5958 22502 6010
rect 22502 5958 22554 6010
rect 22554 5958 22556 6010
rect 22180 5956 22236 5958
rect 22260 5956 22316 5958
rect 22340 5956 22396 5958
rect 22420 5956 22476 5958
rect 22500 5956 22556 5958
rect 24398 15136 24454 15192
rect 28920 30490 28976 30492
rect 29000 30490 29056 30492
rect 29080 30490 29136 30492
rect 29160 30490 29216 30492
rect 29240 30490 29296 30492
rect 28920 30438 28922 30490
rect 28922 30438 28974 30490
rect 28974 30438 28976 30490
rect 29000 30438 29038 30490
rect 29038 30438 29050 30490
rect 29050 30438 29056 30490
rect 29080 30438 29102 30490
rect 29102 30438 29114 30490
rect 29114 30438 29136 30490
rect 29160 30438 29166 30490
rect 29166 30438 29178 30490
rect 29178 30438 29216 30490
rect 29240 30438 29242 30490
rect 29242 30438 29294 30490
rect 29294 30438 29296 30490
rect 28920 30436 28976 30438
rect 29000 30436 29056 30438
rect 29080 30436 29136 30438
rect 29160 30436 29216 30438
rect 29240 30436 29296 30438
rect 28180 29946 28236 29948
rect 28260 29946 28316 29948
rect 28340 29946 28396 29948
rect 28420 29946 28476 29948
rect 28500 29946 28556 29948
rect 28180 29894 28182 29946
rect 28182 29894 28234 29946
rect 28234 29894 28236 29946
rect 28260 29894 28298 29946
rect 28298 29894 28310 29946
rect 28310 29894 28316 29946
rect 28340 29894 28362 29946
rect 28362 29894 28374 29946
rect 28374 29894 28396 29946
rect 28420 29894 28426 29946
rect 28426 29894 28438 29946
rect 28438 29894 28476 29946
rect 28500 29894 28502 29946
rect 28502 29894 28554 29946
rect 28554 29894 28556 29946
rect 28180 29892 28236 29894
rect 28260 29892 28316 29894
rect 28340 29892 28396 29894
rect 28420 29892 28476 29894
rect 28500 29892 28556 29894
rect 28920 29402 28976 29404
rect 29000 29402 29056 29404
rect 29080 29402 29136 29404
rect 29160 29402 29216 29404
rect 29240 29402 29296 29404
rect 28920 29350 28922 29402
rect 28922 29350 28974 29402
rect 28974 29350 28976 29402
rect 29000 29350 29038 29402
rect 29038 29350 29050 29402
rect 29050 29350 29056 29402
rect 29080 29350 29102 29402
rect 29102 29350 29114 29402
rect 29114 29350 29136 29402
rect 29160 29350 29166 29402
rect 29166 29350 29178 29402
rect 29178 29350 29216 29402
rect 29240 29350 29242 29402
rect 29242 29350 29294 29402
rect 29294 29350 29296 29402
rect 28920 29348 28976 29350
rect 29000 29348 29056 29350
rect 29080 29348 29136 29350
rect 29160 29348 29216 29350
rect 29240 29348 29296 29350
rect 28180 28858 28236 28860
rect 28260 28858 28316 28860
rect 28340 28858 28396 28860
rect 28420 28858 28476 28860
rect 28500 28858 28556 28860
rect 28180 28806 28182 28858
rect 28182 28806 28234 28858
rect 28234 28806 28236 28858
rect 28260 28806 28298 28858
rect 28298 28806 28310 28858
rect 28310 28806 28316 28858
rect 28340 28806 28362 28858
rect 28362 28806 28374 28858
rect 28374 28806 28396 28858
rect 28420 28806 28426 28858
rect 28426 28806 28438 28858
rect 28438 28806 28476 28858
rect 28500 28806 28502 28858
rect 28502 28806 28554 28858
rect 28554 28806 28556 28858
rect 28180 28804 28236 28806
rect 28260 28804 28316 28806
rect 28340 28804 28396 28806
rect 28420 28804 28476 28806
rect 28500 28804 28556 28806
rect 28920 28314 28976 28316
rect 29000 28314 29056 28316
rect 29080 28314 29136 28316
rect 29160 28314 29216 28316
rect 29240 28314 29296 28316
rect 28920 28262 28922 28314
rect 28922 28262 28974 28314
rect 28974 28262 28976 28314
rect 29000 28262 29038 28314
rect 29038 28262 29050 28314
rect 29050 28262 29056 28314
rect 29080 28262 29102 28314
rect 29102 28262 29114 28314
rect 29114 28262 29136 28314
rect 29160 28262 29166 28314
rect 29166 28262 29178 28314
rect 29178 28262 29216 28314
rect 29240 28262 29242 28314
rect 29242 28262 29294 28314
rect 29294 28262 29296 28314
rect 28920 28260 28976 28262
rect 29000 28260 29056 28262
rect 29080 28260 29136 28262
rect 29160 28260 29216 28262
rect 29240 28260 29296 28262
rect 28180 27770 28236 27772
rect 28260 27770 28316 27772
rect 28340 27770 28396 27772
rect 28420 27770 28476 27772
rect 28500 27770 28556 27772
rect 28180 27718 28182 27770
rect 28182 27718 28234 27770
rect 28234 27718 28236 27770
rect 28260 27718 28298 27770
rect 28298 27718 28310 27770
rect 28310 27718 28316 27770
rect 28340 27718 28362 27770
rect 28362 27718 28374 27770
rect 28374 27718 28396 27770
rect 28420 27718 28426 27770
rect 28426 27718 28438 27770
rect 28438 27718 28476 27770
rect 28500 27718 28502 27770
rect 28502 27718 28554 27770
rect 28554 27718 28556 27770
rect 28180 27716 28236 27718
rect 28260 27716 28316 27718
rect 28340 27716 28396 27718
rect 28420 27716 28476 27718
rect 28500 27716 28556 27718
rect 22920 5466 22976 5468
rect 23000 5466 23056 5468
rect 23080 5466 23136 5468
rect 23160 5466 23216 5468
rect 23240 5466 23296 5468
rect 22920 5414 22922 5466
rect 22922 5414 22974 5466
rect 22974 5414 22976 5466
rect 23000 5414 23038 5466
rect 23038 5414 23050 5466
rect 23050 5414 23056 5466
rect 23080 5414 23102 5466
rect 23102 5414 23114 5466
rect 23114 5414 23136 5466
rect 23160 5414 23166 5466
rect 23166 5414 23178 5466
rect 23178 5414 23216 5466
rect 23240 5414 23242 5466
rect 23242 5414 23294 5466
rect 23294 5414 23296 5466
rect 22920 5412 22976 5414
rect 23000 5412 23056 5414
rect 23080 5412 23136 5414
rect 23160 5412 23216 5414
rect 23240 5412 23296 5414
rect 25134 8880 25190 8936
rect 22180 4922 22236 4924
rect 22260 4922 22316 4924
rect 22340 4922 22396 4924
rect 22420 4922 22476 4924
rect 22500 4922 22556 4924
rect 22180 4870 22182 4922
rect 22182 4870 22234 4922
rect 22234 4870 22236 4922
rect 22260 4870 22298 4922
rect 22298 4870 22310 4922
rect 22310 4870 22316 4922
rect 22340 4870 22362 4922
rect 22362 4870 22374 4922
rect 22374 4870 22396 4922
rect 22420 4870 22426 4922
rect 22426 4870 22438 4922
rect 22438 4870 22476 4922
rect 22500 4870 22502 4922
rect 22502 4870 22554 4922
rect 22554 4870 22556 4922
rect 22180 4868 22236 4870
rect 22260 4868 22316 4870
rect 22340 4868 22396 4870
rect 22420 4868 22476 4870
rect 22500 4868 22556 4870
rect 22920 4378 22976 4380
rect 23000 4378 23056 4380
rect 23080 4378 23136 4380
rect 23160 4378 23216 4380
rect 23240 4378 23296 4380
rect 22920 4326 22922 4378
rect 22922 4326 22974 4378
rect 22974 4326 22976 4378
rect 23000 4326 23038 4378
rect 23038 4326 23050 4378
rect 23050 4326 23056 4378
rect 23080 4326 23102 4378
rect 23102 4326 23114 4378
rect 23114 4326 23136 4378
rect 23160 4326 23166 4378
rect 23166 4326 23178 4378
rect 23178 4326 23216 4378
rect 23240 4326 23242 4378
rect 23242 4326 23294 4378
rect 23294 4326 23296 4378
rect 22920 4324 22976 4326
rect 23000 4324 23056 4326
rect 23080 4324 23136 4326
rect 23160 4324 23216 4326
rect 23240 4324 23296 4326
rect 28920 27226 28976 27228
rect 29000 27226 29056 27228
rect 29080 27226 29136 27228
rect 29160 27226 29216 27228
rect 29240 27226 29296 27228
rect 28920 27174 28922 27226
rect 28922 27174 28974 27226
rect 28974 27174 28976 27226
rect 29000 27174 29038 27226
rect 29038 27174 29050 27226
rect 29050 27174 29056 27226
rect 29080 27174 29102 27226
rect 29102 27174 29114 27226
rect 29114 27174 29136 27226
rect 29160 27174 29166 27226
rect 29166 27174 29178 27226
rect 29178 27174 29216 27226
rect 29240 27174 29242 27226
rect 29242 27174 29294 27226
rect 29294 27174 29296 27226
rect 28920 27172 28976 27174
rect 29000 27172 29056 27174
rect 29080 27172 29136 27174
rect 29160 27172 29216 27174
rect 29240 27172 29296 27174
rect 28180 26682 28236 26684
rect 28260 26682 28316 26684
rect 28340 26682 28396 26684
rect 28420 26682 28476 26684
rect 28500 26682 28556 26684
rect 28180 26630 28182 26682
rect 28182 26630 28234 26682
rect 28234 26630 28236 26682
rect 28260 26630 28298 26682
rect 28298 26630 28310 26682
rect 28310 26630 28316 26682
rect 28340 26630 28362 26682
rect 28362 26630 28374 26682
rect 28374 26630 28396 26682
rect 28420 26630 28426 26682
rect 28426 26630 28438 26682
rect 28438 26630 28476 26682
rect 28500 26630 28502 26682
rect 28502 26630 28554 26682
rect 28554 26630 28556 26682
rect 28180 26628 28236 26630
rect 28260 26628 28316 26630
rect 28340 26628 28396 26630
rect 28420 26628 28476 26630
rect 28500 26628 28556 26630
rect 28920 26138 28976 26140
rect 29000 26138 29056 26140
rect 29080 26138 29136 26140
rect 29160 26138 29216 26140
rect 29240 26138 29296 26140
rect 28920 26086 28922 26138
rect 28922 26086 28974 26138
rect 28974 26086 28976 26138
rect 29000 26086 29038 26138
rect 29038 26086 29050 26138
rect 29050 26086 29056 26138
rect 29080 26086 29102 26138
rect 29102 26086 29114 26138
rect 29114 26086 29136 26138
rect 29160 26086 29166 26138
rect 29166 26086 29178 26138
rect 29178 26086 29216 26138
rect 29240 26086 29242 26138
rect 29242 26086 29294 26138
rect 29294 26086 29296 26138
rect 28920 26084 28976 26086
rect 29000 26084 29056 26086
rect 29080 26084 29136 26086
rect 29160 26084 29216 26086
rect 29240 26084 29296 26086
rect 28180 25594 28236 25596
rect 28260 25594 28316 25596
rect 28340 25594 28396 25596
rect 28420 25594 28476 25596
rect 28500 25594 28556 25596
rect 28180 25542 28182 25594
rect 28182 25542 28234 25594
rect 28234 25542 28236 25594
rect 28260 25542 28298 25594
rect 28298 25542 28310 25594
rect 28310 25542 28316 25594
rect 28340 25542 28362 25594
rect 28362 25542 28374 25594
rect 28374 25542 28396 25594
rect 28420 25542 28426 25594
rect 28426 25542 28438 25594
rect 28438 25542 28476 25594
rect 28500 25542 28502 25594
rect 28502 25542 28554 25594
rect 28554 25542 28556 25594
rect 28180 25540 28236 25542
rect 28260 25540 28316 25542
rect 28340 25540 28396 25542
rect 28420 25540 28476 25542
rect 28500 25540 28556 25542
rect 28920 25050 28976 25052
rect 29000 25050 29056 25052
rect 29080 25050 29136 25052
rect 29160 25050 29216 25052
rect 29240 25050 29296 25052
rect 28920 24998 28922 25050
rect 28922 24998 28974 25050
rect 28974 24998 28976 25050
rect 29000 24998 29038 25050
rect 29038 24998 29050 25050
rect 29050 24998 29056 25050
rect 29080 24998 29102 25050
rect 29102 24998 29114 25050
rect 29114 24998 29136 25050
rect 29160 24998 29166 25050
rect 29166 24998 29178 25050
rect 29178 24998 29216 25050
rect 29240 24998 29242 25050
rect 29242 24998 29294 25050
rect 29294 24998 29296 25050
rect 28920 24996 28976 24998
rect 29000 24996 29056 24998
rect 29080 24996 29136 24998
rect 29160 24996 29216 24998
rect 29240 24996 29296 24998
rect 28180 24506 28236 24508
rect 28260 24506 28316 24508
rect 28340 24506 28396 24508
rect 28420 24506 28476 24508
rect 28500 24506 28556 24508
rect 28180 24454 28182 24506
rect 28182 24454 28234 24506
rect 28234 24454 28236 24506
rect 28260 24454 28298 24506
rect 28298 24454 28310 24506
rect 28310 24454 28316 24506
rect 28340 24454 28362 24506
rect 28362 24454 28374 24506
rect 28374 24454 28396 24506
rect 28420 24454 28426 24506
rect 28426 24454 28438 24506
rect 28438 24454 28476 24506
rect 28500 24454 28502 24506
rect 28502 24454 28554 24506
rect 28554 24454 28556 24506
rect 28180 24452 28236 24454
rect 28260 24452 28316 24454
rect 28340 24452 28396 24454
rect 28420 24452 28476 24454
rect 28500 24452 28556 24454
rect 28920 23962 28976 23964
rect 29000 23962 29056 23964
rect 29080 23962 29136 23964
rect 29160 23962 29216 23964
rect 29240 23962 29296 23964
rect 28920 23910 28922 23962
rect 28922 23910 28974 23962
rect 28974 23910 28976 23962
rect 29000 23910 29038 23962
rect 29038 23910 29050 23962
rect 29050 23910 29056 23962
rect 29080 23910 29102 23962
rect 29102 23910 29114 23962
rect 29114 23910 29136 23962
rect 29160 23910 29166 23962
rect 29166 23910 29178 23962
rect 29178 23910 29216 23962
rect 29240 23910 29242 23962
rect 29242 23910 29294 23962
rect 29294 23910 29296 23962
rect 28920 23908 28976 23910
rect 29000 23908 29056 23910
rect 29080 23908 29136 23910
rect 29160 23908 29216 23910
rect 29240 23908 29296 23910
rect 28180 23418 28236 23420
rect 28260 23418 28316 23420
rect 28340 23418 28396 23420
rect 28420 23418 28476 23420
rect 28500 23418 28556 23420
rect 28180 23366 28182 23418
rect 28182 23366 28234 23418
rect 28234 23366 28236 23418
rect 28260 23366 28298 23418
rect 28298 23366 28310 23418
rect 28310 23366 28316 23418
rect 28340 23366 28362 23418
rect 28362 23366 28374 23418
rect 28374 23366 28396 23418
rect 28420 23366 28426 23418
rect 28426 23366 28438 23418
rect 28438 23366 28476 23418
rect 28500 23366 28502 23418
rect 28502 23366 28554 23418
rect 28554 23366 28556 23418
rect 28180 23364 28236 23366
rect 28260 23364 28316 23366
rect 28340 23364 28396 23366
rect 28420 23364 28476 23366
rect 28500 23364 28556 23366
rect 28920 22874 28976 22876
rect 29000 22874 29056 22876
rect 29080 22874 29136 22876
rect 29160 22874 29216 22876
rect 29240 22874 29296 22876
rect 28920 22822 28922 22874
rect 28922 22822 28974 22874
rect 28974 22822 28976 22874
rect 29000 22822 29038 22874
rect 29038 22822 29050 22874
rect 29050 22822 29056 22874
rect 29080 22822 29102 22874
rect 29102 22822 29114 22874
rect 29114 22822 29136 22874
rect 29160 22822 29166 22874
rect 29166 22822 29178 22874
rect 29178 22822 29216 22874
rect 29240 22822 29242 22874
rect 29242 22822 29294 22874
rect 29294 22822 29296 22874
rect 28920 22820 28976 22822
rect 29000 22820 29056 22822
rect 29080 22820 29136 22822
rect 29160 22820 29216 22822
rect 29240 22820 29296 22822
rect 28180 22330 28236 22332
rect 28260 22330 28316 22332
rect 28340 22330 28396 22332
rect 28420 22330 28476 22332
rect 28500 22330 28556 22332
rect 28180 22278 28182 22330
rect 28182 22278 28234 22330
rect 28234 22278 28236 22330
rect 28260 22278 28298 22330
rect 28298 22278 28310 22330
rect 28310 22278 28316 22330
rect 28340 22278 28362 22330
rect 28362 22278 28374 22330
rect 28374 22278 28396 22330
rect 28420 22278 28426 22330
rect 28426 22278 28438 22330
rect 28438 22278 28476 22330
rect 28500 22278 28502 22330
rect 28502 22278 28554 22330
rect 28554 22278 28556 22330
rect 28180 22276 28236 22278
rect 28260 22276 28316 22278
rect 28340 22276 28396 22278
rect 28420 22276 28476 22278
rect 28500 22276 28556 22278
rect 28920 21786 28976 21788
rect 29000 21786 29056 21788
rect 29080 21786 29136 21788
rect 29160 21786 29216 21788
rect 29240 21786 29296 21788
rect 28920 21734 28922 21786
rect 28922 21734 28974 21786
rect 28974 21734 28976 21786
rect 29000 21734 29038 21786
rect 29038 21734 29050 21786
rect 29050 21734 29056 21786
rect 29080 21734 29102 21786
rect 29102 21734 29114 21786
rect 29114 21734 29136 21786
rect 29160 21734 29166 21786
rect 29166 21734 29178 21786
rect 29178 21734 29216 21786
rect 29240 21734 29242 21786
rect 29242 21734 29294 21786
rect 29294 21734 29296 21786
rect 28920 21732 28976 21734
rect 29000 21732 29056 21734
rect 29080 21732 29136 21734
rect 29160 21732 29216 21734
rect 29240 21732 29296 21734
rect 28180 21242 28236 21244
rect 28260 21242 28316 21244
rect 28340 21242 28396 21244
rect 28420 21242 28476 21244
rect 28500 21242 28556 21244
rect 28180 21190 28182 21242
rect 28182 21190 28234 21242
rect 28234 21190 28236 21242
rect 28260 21190 28298 21242
rect 28298 21190 28310 21242
rect 28310 21190 28316 21242
rect 28340 21190 28362 21242
rect 28362 21190 28374 21242
rect 28374 21190 28396 21242
rect 28420 21190 28426 21242
rect 28426 21190 28438 21242
rect 28438 21190 28476 21242
rect 28500 21190 28502 21242
rect 28502 21190 28554 21242
rect 28554 21190 28556 21242
rect 28180 21188 28236 21190
rect 28260 21188 28316 21190
rect 28340 21188 28396 21190
rect 28420 21188 28476 21190
rect 28500 21188 28556 21190
rect 28920 20698 28976 20700
rect 29000 20698 29056 20700
rect 29080 20698 29136 20700
rect 29160 20698 29216 20700
rect 29240 20698 29296 20700
rect 28920 20646 28922 20698
rect 28922 20646 28974 20698
rect 28974 20646 28976 20698
rect 29000 20646 29038 20698
rect 29038 20646 29050 20698
rect 29050 20646 29056 20698
rect 29080 20646 29102 20698
rect 29102 20646 29114 20698
rect 29114 20646 29136 20698
rect 29160 20646 29166 20698
rect 29166 20646 29178 20698
rect 29178 20646 29216 20698
rect 29240 20646 29242 20698
rect 29242 20646 29294 20698
rect 29294 20646 29296 20698
rect 28920 20644 28976 20646
rect 29000 20644 29056 20646
rect 29080 20644 29136 20646
rect 29160 20644 29216 20646
rect 29240 20644 29296 20646
rect 28180 20154 28236 20156
rect 28260 20154 28316 20156
rect 28340 20154 28396 20156
rect 28420 20154 28476 20156
rect 28500 20154 28556 20156
rect 28180 20102 28182 20154
rect 28182 20102 28234 20154
rect 28234 20102 28236 20154
rect 28260 20102 28298 20154
rect 28298 20102 28310 20154
rect 28310 20102 28316 20154
rect 28340 20102 28362 20154
rect 28362 20102 28374 20154
rect 28374 20102 28396 20154
rect 28420 20102 28426 20154
rect 28426 20102 28438 20154
rect 28438 20102 28476 20154
rect 28500 20102 28502 20154
rect 28502 20102 28554 20154
rect 28554 20102 28556 20154
rect 28180 20100 28236 20102
rect 28260 20100 28316 20102
rect 28340 20100 28396 20102
rect 28420 20100 28476 20102
rect 28500 20100 28556 20102
rect 28920 19610 28976 19612
rect 29000 19610 29056 19612
rect 29080 19610 29136 19612
rect 29160 19610 29216 19612
rect 29240 19610 29296 19612
rect 28920 19558 28922 19610
rect 28922 19558 28974 19610
rect 28974 19558 28976 19610
rect 29000 19558 29038 19610
rect 29038 19558 29050 19610
rect 29050 19558 29056 19610
rect 29080 19558 29102 19610
rect 29102 19558 29114 19610
rect 29114 19558 29136 19610
rect 29160 19558 29166 19610
rect 29166 19558 29178 19610
rect 29178 19558 29216 19610
rect 29240 19558 29242 19610
rect 29242 19558 29294 19610
rect 29294 19558 29296 19610
rect 28920 19556 28976 19558
rect 29000 19556 29056 19558
rect 29080 19556 29136 19558
rect 29160 19556 29216 19558
rect 29240 19556 29296 19558
rect 28180 19066 28236 19068
rect 28260 19066 28316 19068
rect 28340 19066 28396 19068
rect 28420 19066 28476 19068
rect 28500 19066 28556 19068
rect 28180 19014 28182 19066
rect 28182 19014 28234 19066
rect 28234 19014 28236 19066
rect 28260 19014 28298 19066
rect 28298 19014 28310 19066
rect 28310 19014 28316 19066
rect 28340 19014 28362 19066
rect 28362 19014 28374 19066
rect 28374 19014 28396 19066
rect 28420 19014 28426 19066
rect 28426 19014 28438 19066
rect 28438 19014 28476 19066
rect 28500 19014 28502 19066
rect 28502 19014 28554 19066
rect 28554 19014 28556 19066
rect 28180 19012 28236 19014
rect 28260 19012 28316 19014
rect 28340 19012 28396 19014
rect 28420 19012 28476 19014
rect 28500 19012 28556 19014
rect 28920 18522 28976 18524
rect 29000 18522 29056 18524
rect 29080 18522 29136 18524
rect 29160 18522 29216 18524
rect 29240 18522 29296 18524
rect 28920 18470 28922 18522
rect 28922 18470 28974 18522
rect 28974 18470 28976 18522
rect 29000 18470 29038 18522
rect 29038 18470 29050 18522
rect 29050 18470 29056 18522
rect 29080 18470 29102 18522
rect 29102 18470 29114 18522
rect 29114 18470 29136 18522
rect 29160 18470 29166 18522
rect 29166 18470 29178 18522
rect 29178 18470 29216 18522
rect 29240 18470 29242 18522
rect 29242 18470 29294 18522
rect 29294 18470 29296 18522
rect 28920 18468 28976 18470
rect 29000 18468 29056 18470
rect 29080 18468 29136 18470
rect 29160 18468 29216 18470
rect 29240 18468 29296 18470
rect 28180 17978 28236 17980
rect 28260 17978 28316 17980
rect 28340 17978 28396 17980
rect 28420 17978 28476 17980
rect 28500 17978 28556 17980
rect 28180 17926 28182 17978
rect 28182 17926 28234 17978
rect 28234 17926 28236 17978
rect 28260 17926 28298 17978
rect 28298 17926 28310 17978
rect 28310 17926 28316 17978
rect 28340 17926 28362 17978
rect 28362 17926 28374 17978
rect 28374 17926 28396 17978
rect 28420 17926 28426 17978
rect 28426 17926 28438 17978
rect 28438 17926 28476 17978
rect 28500 17926 28502 17978
rect 28502 17926 28554 17978
rect 28554 17926 28556 17978
rect 28180 17924 28236 17926
rect 28260 17924 28316 17926
rect 28340 17924 28396 17926
rect 28420 17924 28476 17926
rect 28500 17924 28556 17926
rect 28920 17434 28976 17436
rect 29000 17434 29056 17436
rect 29080 17434 29136 17436
rect 29160 17434 29216 17436
rect 29240 17434 29296 17436
rect 28920 17382 28922 17434
rect 28922 17382 28974 17434
rect 28974 17382 28976 17434
rect 29000 17382 29038 17434
rect 29038 17382 29050 17434
rect 29050 17382 29056 17434
rect 29080 17382 29102 17434
rect 29102 17382 29114 17434
rect 29114 17382 29136 17434
rect 29160 17382 29166 17434
rect 29166 17382 29178 17434
rect 29178 17382 29216 17434
rect 29240 17382 29242 17434
rect 29242 17382 29294 17434
rect 29294 17382 29296 17434
rect 28920 17380 28976 17382
rect 29000 17380 29056 17382
rect 29080 17380 29136 17382
rect 29160 17380 29216 17382
rect 29240 17380 29296 17382
rect 28180 16890 28236 16892
rect 28260 16890 28316 16892
rect 28340 16890 28396 16892
rect 28420 16890 28476 16892
rect 28500 16890 28556 16892
rect 28180 16838 28182 16890
rect 28182 16838 28234 16890
rect 28234 16838 28236 16890
rect 28260 16838 28298 16890
rect 28298 16838 28310 16890
rect 28310 16838 28316 16890
rect 28340 16838 28362 16890
rect 28362 16838 28374 16890
rect 28374 16838 28396 16890
rect 28420 16838 28426 16890
rect 28426 16838 28438 16890
rect 28438 16838 28476 16890
rect 28500 16838 28502 16890
rect 28502 16838 28554 16890
rect 28554 16838 28556 16890
rect 28180 16836 28236 16838
rect 28260 16836 28316 16838
rect 28340 16836 28396 16838
rect 28420 16836 28476 16838
rect 28500 16836 28556 16838
rect 28920 16346 28976 16348
rect 29000 16346 29056 16348
rect 29080 16346 29136 16348
rect 29160 16346 29216 16348
rect 29240 16346 29296 16348
rect 28920 16294 28922 16346
rect 28922 16294 28974 16346
rect 28974 16294 28976 16346
rect 29000 16294 29038 16346
rect 29038 16294 29050 16346
rect 29050 16294 29056 16346
rect 29080 16294 29102 16346
rect 29102 16294 29114 16346
rect 29114 16294 29136 16346
rect 29160 16294 29166 16346
rect 29166 16294 29178 16346
rect 29178 16294 29216 16346
rect 29240 16294 29242 16346
rect 29242 16294 29294 16346
rect 29294 16294 29296 16346
rect 28920 16292 28976 16294
rect 29000 16292 29056 16294
rect 29080 16292 29136 16294
rect 29160 16292 29216 16294
rect 29240 16292 29296 16294
rect 28180 15802 28236 15804
rect 28260 15802 28316 15804
rect 28340 15802 28396 15804
rect 28420 15802 28476 15804
rect 28500 15802 28556 15804
rect 28180 15750 28182 15802
rect 28182 15750 28234 15802
rect 28234 15750 28236 15802
rect 28260 15750 28298 15802
rect 28298 15750 28310 15802
rect 28310 15750 28316 15802
rect 28340 15750 28362 15802
rect 28362 15750 28374 15802
rect 28374 15750 28396 15802
rect 28420 15750 28426 15802
rect 28426 15750 28438 15802
rect 28438 15750 28476 15802
rect 28500 15750 28502 15802
rect 28502 15750 28554 15802
rect 28554 15750 28556 15802
rect 28180 15748 28236 15750
rect 28260 15748 28316 15750
rect 28340 15748 28396 15750
rect 28420 15748 28476 15750
rect 28500 15748 28556 15750
rect 28920 15258 28976 15260
rect 29000 15258 29056 15260
rect 29080 15258 29136 15260
rect 29160 15258 29216 15260
rect 29240 15258 29296 15260
rect 28920 15206 28922 15258
rect 28922 15206 28974 15258
rect 28974 15206 28976 15258
rect 29000 15206 29038 15258
rect 29038 15206 29050 15258
rect 29050 15206 29056 15258
rect 29080 15206 29102 15258
rect 29102 15206 29114 15258
rect 29114 15206 29136 15258
rect 29160 15206 29166 15258
rect 29166 15206 29178 15258
rect 29178 15206 29216 15258
rect 29240 15206 29242 15258
rect 29242 15206 29294 15258
rect 29294 15206 29296 15258
rect 28920 15204 28976 15206
rect 29000 15204 29056 15206
rect 29080 15204 29136 15206
rect 29160 15204 29216 15206
rect 29240 15204 29296 15206
rect 28180 14714 28236 14716
rect 28260 14714 28316 14716
rect 28340 14714 28396 14716
rect 28420 14714 28476 14716
rect 28500 14714 28556 14716
rect 28180 14662 28182 14714
rect 28182 14662 28234 14714
rect 28234 14662 28236 14714
rect 28260 14662 28298 14714
rect 28298 14662 28310 14714
rect 28310 14662 28316 14714
rect 28340 14662 28362 14714
rect 28362 14662 28374 14714
rect 28374 14662 28396 14714
rect 28420 14662 28426 14714
rect 28426 14662 28438 14714
rect 28438 14662 28476 14714
rect 28500 14662 28502 14714
rect 28502 14662 28554 14714
rect 28554 14662 28556 14714
rect 28180 14660 28236 14662
rect 28260 14660 28316 14662
rect 28340 14660 28396 14662
rect 28420 14660 28476 14662
rect 28500 14660 28556 14662
rect 28920 14170 28976 14172
rect 29000 14170 29056 14172
rect 29080 14170 29136 14172
rect 29160 14170 29216 14172
rect 29240 14170 29296 14172
rect 28920 14118 28922 14170
rect 28922 14118 28974 14170
rect 28974 14118 28976 14170
rect 29000 14118 29038 14170
rect 29038 14118 29050 14170
rect 29050 14118 29056 14170
rect 29080 14118 29102 14170
rect 29102 14118 29114 14170
rect 29114 14118 29136 14170
rect 29160 14118 29166 14170
rect 29166 14118 29178 14170
rect 29178 14118 29216 14170
rect 29240 14118 29242 14170
rect 29242 14118 29294 14170
rect 29294 14118 29296 14170
rect 28920 14116 28976 14118
rect 29000 14116 29056 14118
rect 29080 14116 29136 14118
rect 29160 14116 29216 14118
rect 29240 14116 29296 14118
rect 28180 13626 28236 13628
rect 28260 13626 28316 13628
rect 28340 13626 28396 13628
rect 28420 13626 28476 13628
rect 28500 13626 28556 13628
rect 28180 13574 28182 13626
rect 28182 13574 28234 13626
rect 28234 13574 28236 13626
rect 28260 13574 28298 13626
rect 28298 13574 28310 13626
rect 28310 13574 28316 13626
rect 28340 13574 28362 13626
rect 28362 13574 28374 13626
rect 28374 13574 28396 13626
rect 28420 13574 28426 13626
rect 28426 13574 28438 13626
rect 28438 13574 28476 13626
rect 28500 13574 28502 13626
rect 28502 13574 28554 13626
rect 28554 13574 28556 13626
rect 28180 13572 28236 13574
rect 28260 13572 28316 13574
rect 28340 13572 28396 13574
rect 28420 13572 28476 13574
rect 28500 13572 28556 13574
rect 28920 13082 28976 13084
rect 29000 13082 29056 13084
rect 29080 13082 29136 13084
rect 29160 13082 29216 13084
rect 29240 13082 29296 13084
rect 28920 13030 28922 13082
rect 28922 13030 28974 13082
rect 28974 13030 28976 13082
rect 29000 13030 29038 13082
rect 29038 13030 29050 13082
rect 29050 13030 29056 13082
rect 29080 13030 29102 13082
rect 29102 13030 29114 13082
rect 29114 13030 29136 13082
rect 29160 13030 29166 13082
rect 29166 13030 29178 13082
rect 29178 13030 29216 13082
rect 29240 13030 29242 13082
rect 29242 13030 29294 13082
rect 29294 13030 29296 13082
rect 28920 13028 28976 13030
rect 29000 13028 29056 13030
rect 29080 13028 29136 13030
rect 29160 13028 29216 13030
rect 29240 13028 29296 13030
rect 28180 12538 28236 12540
rect 28260 12538 28316 12540
rect 28340 12538 28396 12540
rect 28420 12538 28476 12540
rect 28500 12538 28556 12540
rect 28180 12486 28182 12538
rect 28182 12486 28234 12538
rect 28234 12486 28236 12538
rect 28260 12486 28298 12538
rect 28298 12486 28310 12538
rect 28310 12486 28316 12538
rect 28340 12486 28362 12538
rect 28362 12486 28374 12538
rect 28374 12486 28396 12538
rect 28420 12486 28426 12538
rect 28426 12486 28438 12538
rect 28438 12486 28476 12538
rect 28500 12486 28502 12538
rect 28502 12486 28554 12538
rect 28554 12486 28556 12538
rect 28180 12484 28236 12486
rect 28260 12484 28316 12486
rect 28340 12484 28396 12486
rect 28420 12484 28476 12486
rect 28500 12484 28556 12486
rect 31298 25200 31354 25256
rect 30930 19116 30932 19136
rect 30932 19116 30984 19136
rect 30984 19116 30986 19136
rect 30930 19080 30986 19116
rect 31298 12960 31354 13016
rect 28920 11994 28976 11996
rect 29000 11994 29056 11996
rect 29080 11994 29136 11996
rect 29160 11994 29216 11996
rect 29240 11994 29296 11996
rect 28920 11942 28922 11994
rect 28922 11942 28974 11994
rect 28974 11942 28976 11994
rect 29000 11942 29038 11994
rect 29038 11942 29050 11994
rect 29050 11942 29056 11994
rect 29080 11942 29102 11994
rect 29102 11942 29114 11994
rect 29114 11942 29136 11994
rect 29160 11942 29166 11994
rect 29166 11942 29178 11994
rect 29178 11942 29216 11994
rect 29240 11942 29242 11994
rect 29242 11942 29294 11994
rect 29294 11942 29296 11994
rect 28920 11940 28976 11942
rect 29000 11940 29056 11942
rect 29080 11940 29136 11942
rect 29160 11940 29216 11942
rect 29240 11940 29296 11942
rect 28180 11450 28236 11452
rect 28260 11450 28316 11452
rect 28340 11450 28396 11452
rect 28420 11450 28476 11452
rect 28500 11450 28556 11452
rect 28180 11398 28182 11450
rect 28182 11398 28234 11450
rect 28234 11398 28236 11450
rect 28260 11398 28298 11450
rect 28298 11398 28310 11450
rect 28310 11398 28316 11450
rect 28340 11398 28362 11450
rect 28362 11398 28374 11450
rect 28374 11398 28396 11450
rect 28420 11398 28426 11450
rect 28426 11398 28438 11450
rect 28438 11398 28476 11450
rect 28500 11398 28502 11450
rect 28502 11398 28554 11450
rect 28554 11398 28556 11450
rect 28180 11396 28236 11398
rect 28260 11396 28316 11398
rect 28340 11396 28396 11398
rect 28420 11396 28476 11398
rect 28500 11396 28556 11398
rect 28920 10906 28976 10908
rect 29000 10906 29056 10908
rect 29080 10906 29136 10908
rect 29160 10906 29216 10908
rect 29240 10906 29296 10908
rect 28920 10854 28922 10906
rect 28922 10854 28974 10906
rect 28974 10854 28976 10906
rect 29000 10854 29038 10906
rect 29038 10854 29050 10906
rect 29050 10854 29056 10906
rect 29080 10854 29102 10906
rect 29102 10854 29114 10906
rect 29114 10854 29136 10906
rect 29160 10854 29166 10906
rect 29166 10854 29178 10906
rect 29178 10854 29216 10906
rect 29240 10854 29242 10906
rect 29242 10854 29294 10906
rect 29294 10854 29296 10906
rect 28920 10852 28976 10854
rect 29000 10852 29056 10854
rect 29080 10852 29136 10854
rect 29160 10852 29216 10854
rect 29240 10852 29296 10854
rect 28180 10362 28236 10364
rect 28260 10362 28316 10364
rect 28340 10362 28396 10364
rect 28420 10362 28476 10364
rect 28500 10362 28556 10364
rect 28180 10310 28182 10362
rect 28182 10310 28234 10362
rect 28234 10310 28236 10362
rect 28260 10310 28298 10362
rect 28298 10310 28310 10362
rect 28310 10310 28316 10362
rect 28340 10310 28362 10362
rect 28362 10310 28374 10362
rect 28374 10310 28396 10362
rect 28420 10310 28426 10362
rect 28426 10310 28438 10362
rect 28438 10310 28476 10362
rect 28500 10310 28502 10362
rect 28502 10310 28554 10362
rect 28554 10310 28556 10362
rect 28180 10308 28236 10310
rect 28260 10308 28316 10310
rect 28340 10308 28396 10310
rect 28420 10308 28476 10310
rect 28500 10308 28556 10310
rect 28920 9818 28976 9820
rect 29000 9818 29056 9820
rect 29080 9818 29136 9820
rect 29160 9818 29216 9820
rect 29240 9818 29296 9820
rect 28920 9766 28922 9818
rect 28922 9766 28974 9818
rect 28974 9766 28976 9818
rect 29000 9766 29038 9818
rect 29038 9766 29050 9818
rect 29050 9766 29056 9818
rect 29080 9766 29102 9818
rect 29102 9766 29114 9818
rect 29114 9766 29136 9818
rect 29160 9766 29166 9818
rect 29166 9766 29178 9818
rect 29178 9766 29216 9818
rect 29240 9766 29242 9818
rect 29242 9766 29294 9818
rect 29294 9766 29296 9818
rect 28920 9764 28976 9766
rect 29000 9764 29056 9766
rect 29080 9764 29136 9766
rect 29160 9764 29216 9766
rect 29240 9764 29296 9766
rect 28180 9274 28236 9276
rect 28260 9274 28316 9276
rect 28340 9274 28396 9276
rect 28420 9274 28476 9276
rect 28500 9274 28556 9276
rect 28180 9222 28182 9274
rect 28182 9222 28234 9274
rect 28234 9222 28236 9274
rect 28260 9222 28298 9274
rect 28298 9222 28310 9274
rect 28310 9222 28316 9274
rect 28340 9222 28362 9274
rect 28362 9222 28374 9274
rect 28374 9222 28396 9274
rect 28420 9222 28426 9274
rect 28426 9222 28438 9274
rect 28438 9222 28476 9274
rect 28500 9222 28502 9274
rect 28502 9222 28554 9274
rect 28554 9222 28556 9274
rect 28180 9220 28236 9222
rect 28260 9220 28316 9222
rect 28340 9220 28396 9222
rect 28420 9220 28476 9222
rect 28500 9220 28556 9222
rect 28920 8730 28976 8732
rect 29000 8730 29056 8732
rect 29080 8730 29136 8732
rect 29160 8730 29216 8732
rect 29240 8730 29296 8732
rect 28920 8678 28922 8730
rect 28922 8678 28974 8730
rect 28974 8678 28976 8730
rect 29000 8678 29038 8730
rect 29038 8678 29050 8730
rect 29050 8678 29056 8730
rect 29080 8678 29102 8730
rect 29102 8678 29114 8730
rect 29114 8678 29136 8730
rect 29160 8678 29166 8730
rect 29166 8678 29178 8730
rect 29178 8678 29216 8730
rect 29240 8678 29242 8730
rect 29242 8678 29294 8730
rect 29294 8678 29296 8730
rect 28920 8676 28976 8678
rect 29000 8676 29056 8678
rect 29080 8676 29136 8678
rect 29160 8676 29216 8678
rect 29240 8676 29296 8678
rect 28180 8186 28236 8188
rect 28260 8186 28316 8188
rect 28340 8186 28396 8188
rect 28420 8186 28476 8188
rect 28500 8186 28556 8188
rect 28180 8134 28182 8186
rect 28182 8134 28234 8186
rect 28234 8134 28236 8186
rect 28260 8134 28298 8186
rect 28298 8134 28310 8186
rect 28310 8134 28316 8186
rect 28340 8134 28362 8186
rect 28362 8134 28374 8186
rect 28374 8134 28396 8186
rect 28420 8134 28426 8186
rect 28426 8134 28438 8186
rect 28438 8134 28476 8186
rect 28500 8134 28502 8186
rect 28502 8134 28554 8186
rect 28554 8134 28556 8186
rect 28180 8132 28236 8134
rect 28260 8132 28316 8134
rect 28340 8132 28396 8134
rect 28420 8132 28476 8134
rect 28500 8132 28556 8134
rect 28920 7642 28976 7644
rect 29000 7642 29056 7644
rect 29080 7642 29136 7644
rect 29160 7642 29216 7644
rect 29240 7642 29296 7644
rect 28920 7590 28922 7642
rect 28922 7590 28974 7642
rect 28974 7590 28976 7642
rect 29000 7590 29038 7642
rect 29038 7590 29050 7642
rect 29050 7590 29056 7642
rect 29080 7590 29102 7642
rect 29102 7590 29114 7642
rect 29114 7590 29136 7642
rect 29160 7590 29166 7642
rect 29166 7590 29178 7642
rect 29178 7590 29216 7642
rect 29240 7590 29242 7642
rect 29242 7590 29294 7642
rect 29294 7590 29296 7642
rect 28920 7588 28976 7590
rect 29000 7588 29056 7590
rect 29080 7588 29136 7590
rect 29160 7588 29216 7590
rect 29240 7588 29296 7590
rect 31298 7520 31354 7576
rect 28180 7098 28236 7100
rect 28260 7098 28316 7100
rect 28340 7098 28396 7100
rect 28420 7098 28476 7100
rect 28500 7098 28556 7100
rect 28180 7046 28182 7098
rect 28182 7046 28234 7098
rect 28234 7046 28236 7098
rect 28260 7046 28298 7098
rect 28298 7046 28310 7098
rect 28310 7046 28316 7098
rect 28340 7046 28362 7098
rect 28362 7046 28374 7098
rect 28374 7046 28396 7098
rect 28420 7046 28426 7098
rect 28426 7046 28438 7098
rect 28438 7046 28476 7098
rect 28500 7046 28502 7098
rect 28502 7046 28554 7098
rect 28554 7046 28556 7098
rect 28180 7044 28236 7046
rect 28260 7044 28316 7046
rect 28340 7044 28396 7046
rect 28420 7044 28476 7046
rect 28500 7044 28556 7046
rect 28920 6554 28976 6556
rect 29000 6554 29056 6556
rect 29080 6554 29136 6556
rect 29160 6554 29216 6556
rect 29240 6554 29296 6556
rect 28920 6502 28922 6554
rect 28922 6502 28974 6554
rect 28974 6502 28976 6554
rect 29000 6502 29038 6554
rect 29038 6502 29050 6554
rect 29050 6502 29056 6554
rect 29080 6502 29102 6554
rect 29102 6502 29114 6554
rect 29114 6502 29136 6554
rect 29160 6502 29166 6554
rect 29166 6502 29178 6554
rect 29178 6502 29216 6554
rect 29240 6502 29242 6554
rect 29242 6502 29294 6554
rect 29294 6502 29296 6554
rect 28920 6500 28976 6502
rect 29000 6500 29056 6502
rect 29080 6500 29136 6502
rect 29160 6500 29216 6502
rect 29240 6500 29296 6502
rect 28180 6010 28236 6012
rect 28260 6010 28316 6012
rect 28340 6010 28396 6012
rect 28420 6010 28476 6012
rect 28500 6010 28556 6012
rect 28180 5958 28182 6010
rect 28182 5958 28234 6010
rect 28234 5958 28236 6010
rect 28260 5958 28298 6010
rect 28298 5958 28310 6010
rect 28310 5958 28316 6010
rect 28340 5958 28362 6010
rect 28362 5958 28374 6010
rect 28374 5958 28396 6010
rect 28420 5958 28426 6010
rect 28426 5958 28438 6010
rect 28438 5958 28476 6010
rect 28500 5958 28502 6010
rect 28502 5958 28554 6010
rect 28554 5958 28556 6010
rect 28180 5956 28236 5958
rect 28260 5956 28316 5958
rect 28340 5956 28396 5958
rect 28420 5956 28476 5958
rect 28500 5956 28556 5958
rect 28920 5466 28976 5468
rect 29000 5466 29056 5468
rect 29080 5466 29136 5468
rect 29160 5466 29216 5468
rect 29240 5466 29296 5468
rect 28920 5414 28922 5466
rect 28922 5414 28974 5466
rect 28974 5414 28976 5466
rect 29000 5414 29038 5466
rect 29038 5414 29050 5466
rect 29050 5414 29056 5466
rect 29080 5414 29102 5466
rect 29102 5414 29114 5466
rect 29114 5414 29136 5466
rect 29160 5414 29166 5466
rect 29166 5414 29178 5466
rect 29178 5414 29216 5466
rect 29240 5414 29242 5466
rect 29242 5414 29294 5466
rect 29294 5414 29296 5466
rect 28920 5412 28976 5414
rect 29000 5412 29056 5414
rect 29080 5412 29136 5414
rect 29160 5412 29216 5414
rect 29240 5412 29296 5414
rect 22180 3834 22236 3836
rect 22260 3834 22316 3836
rect 22340 3834 22396 3836
rect 22420 3834 22476 3836
rect 22500 3834 22556 3836
rect 22180 3782 22182 3834
rect 22182 3782 22234 3834
rect 22234 3782 22236 3834
rect 22260 3782 22298 3834
rect 22298 3782 22310 3834
rect 22310 3782 22316 3834
rect 22340 3782 22362 3834
rect 22362 3782 22374 3834
rect 22374 3782 22396 3834
rect 22420 3782 22426 3834
rect 22426 3782 22438 3834
rect 22438 3782 22476 3834
rect 22500 3782 22502 3834
rect 22502 3782 22554 3834
rect 22554 3782 22556 3834
rect 22180 3780 22236 3782
rect 22260 3780 22316 3782
rect 22340 3780 22396 3782
rect 22420 3780 22476 3782
rect 22500 3780 22556 3782
rect 28180 4922 28236 4924
rect 28260 4922 28316 4924
rect 28340 4922 28396 4924
rect 28420 4922 28476 4924
rect 28500 4922 28556 4924
rect 28180 4870 28182 4922
rect 28182 4870 28234 4922
rect 28234 4870 28236 4922
rect 28260 4870 28298 4922
rect 28298 4870 28310 4922
rect 28310 4870 28316 4922
rect 28340 4870 28362 4922
rect 28362 4870 28374 4922
rect 28374 4870 28396 4922
rect 28420 4870 28426 4922
rect 28426 4870 28438 4922
rect 28438 4870 28476 4922
rect 28500 4870 28502 4922
rect 28502 4870 28554 4922
rect 28554 4870 28556 4922
rect 28180 4868 28236 4870
rect 28260 4868 28316 4870
rect 28340 4868 28396 4870
rect 28420 4868 28476 4870
rect 28500 4868 28556 4870
rect 28920 4378 28976 4380
rect 29000 4378 29056 4380
rect 29080 4378 29136 4380
rect 29160 4378 29216 4380
rect 29240 4378 29296 4380
rect 28920 4326 28922 4378
rect 28922 4326 28974 4378
rect 28974 4326 28976 4378
rect 29000 4326 29038 4378
rect 29038 4326 29050 4378
rect 29050 4326 29056 4378
rect 29080 4326 29102 4378
rect 29102 4326 29114 4378
rect 29114 4326 29136 4378
rect 29160 4326 29166 4378
rect 29166 4326 29178 4378
rect 29178 4326 29216 4378
rect 29240 4326 29242 4378
rect 29242 4326 29294 4378
rect 29294 4326 29296 4378
rect 28920 4324 28976 4326
rect 29000 4324 29056 4326
rect 29080 4324 29136 4326
rect 29160 4324 29216 4326
rect 29240 4324 29296 4326
rect 28180 3834 28236 3836
rect 28260 3834 28316 3836
rect 28340 3834 28396 3836
rect 28420 3834 28476 3836
rect 28500 3834 28556 3836
rect 28180 3782 28182 3834
rect 28182 3782 28234 3834
rect 28234 3782 28236 3834
rect 28260 3782 28298 3834
rect 28298 3782 28310 3834
rect 28310 3782 28316 3834
rect 28340 3782 28362 3834
rect 28362 3782 28374 3834
rect 28374 3782 28396 3834
rect 28420 3782 28426 3834
rect 28426 3782 28438 3834
rect 28438 3782 28476 3834
rect 28500 3782 28502 3834
rect 28502 3782 28554 3834
rect 28554 3782 28556 3834
rect 28180 3780 28236 3782
rect 28260 3780 28316 3782
rect 28340 3780 28396 3782
rect 28420 3780 28476 3782
rect 28500 3780 28556 3782
rect 16180 2746 16236 2748
rect 16260 2746 16316 2748
rect 16340 2746 16396 2748
rect 16420 2746 16476 2748
rect 16500 2746 16556 2748
rect 16180 2694 16182 2746
rect 16182 2694 16234 2746
rect 16234 2694 16236 2746
rect 16260 2694 16298 2746
rect 16298 2694 16310 2746
rect 16310 2694 16316 2746
rect 16340 2694 16362 2746
rect 16362 2694 16374 2746
rect 16374 2694 16396 2746
rect 16420 2694 16426 2746
rect 16426 2694 16438 2746
rect 16438 2694 16476 2746
rect 16500 2694 16502 2746
rect 16502 2694 16554 2746
rect 16554 2694 16556 2746
rect 16180 2692 16236 2694
rect 16260 2692 16316 2694
rect 16340 2692 16396 2694
rect 16420 2692 16476 2694
rect 16500 2692 16556 2694
rect 22920 3290 22976 3292
rect 23000 3290 23056 3292
rect 23080 3290 23136 3292
rect 23160 3290 23216 3292
rect 23240 3290 23296 3292
rect 22920 3238 22922 3290
rect 22922 3238 22974 3290
rect 22974 3238 22976 3290
rect 23000 3238 23038 3290
rect 23038 3238 23050 3290
rect 23050 3238 23056 3290
rect 23080 3238 23102 3290
rect 23102 3238 23114 3290
rect 23114 3238 23136 3290
rect 23160 3238 23166 3290
rect 23166 3238 23178 3290
rect 23178 3238 23216 3290
rect 23240 3238 23242 3290
rect 23242 3238 23294 3290
rect 23294 3238 23296 3290
rect 22920 3236 22976 3238
rect 23000 3236 23056 3238
rect 23080 3236 23136 3238
rect 23160 3236 23216 3238
rect 23240 3236 23296 3238
rect 22180 2746 22236 2748
rect 22260 2746 22316 2748
rect 22340 2746 22396 2748
rect 22420 2746 22476 2748
rect 22500 2746 22556 2748
rect 22180 2694 22182 2746
rect 22182 2694 22234 2746
rect 22234 2694 22236 2746
rect 22260 2694 22298 2746
rect 22298 2694 22310 2746
rect 22310 2694 22316 2746
rect 22340 2694 22362 2746
rect 22362 2694 22374 2746
rect 22374 2694 22396 2746
rect 22420 2694 22426 2746
rect 22426 2694 22438 2746
rect 22438 2694 22476 2746
rect 22500 2694 22502 2746
rect 22502 2694 22554 2746
rect 22554 2694 22556 2746
rect 22180 2692 22236 2694
rect 22260 2692 22316 2694
rect 22340 2692 22396 2694
rect 22420 2692 22476 2694
rect 22500 2692 22556 2694
rect 28180 2746 28236 2748
rect 28260 2746 28316 2748
rect 28340 2746 28396 2748
rect 28420 2746 28476 2748
rect 28500 2746 28556 2748
rect 28180 2694 28182 2746
rect 28182 2694 28234 2746
rect 28234 2694 28236 2746
rect 28260 2694 28298 2746
rect 28298 2694 28310 2746
rect 28310 2694 28316 2746
rect 28340 2694 28362 2746
rect 28362 2694 28374 2746
rect 28374 2694 28396 2746
rect 28420 2694 28426 2746
rect 28426 2694 28438 2746
rect 28438 2694 28476 2746
rect 28500 2694 28502 2746
rect 28502 2694 28554 2746
rect 28554 2694 28556 2746
rect 28180 2692 28236 2694
rect 28260 2692 28316 2694
rect 28340 2692 28396 2694
rect 28420 2692 28476 2694
rect 28500 2692 28556 2694
rect 28920 3290 28976 3292
rect 29000 3290 29056 3292
rect 29080 3290 29136 3292
rect 29160 3290 29216 3292
rect 29240 3290 29296 3292
rect 28920 3238 28922 3290
rect 28922 3238 28974 3290
rect 28974 3238 28976 3290
rect 29000 3238 29038 3290
rect 29038 3238 29050 3290
rect 29050 3238 29056 3290
rect 29080 3238 29102 3290
rect 29102 3238 29114 3290
rect 29114 3238 29136 3290
rect 29160 3238 29166 3290
rect 29166 3238 29178 3290
rect 29178 3238 29216 3290
rect 29240 3238 29242 3290
rect 29242 3238 29294 3290
rect 29294 3238 29296 3290
rect 28920 3236 28976 3238
rect 29000 3236 29056 3238
rect 29080 3236 29136 3238
rect 29160 3236 29216 3238
rect 29240 3236 29296 3238
rect 4920 2202 4976 2204
rect 5000 2202 5056 2204
rect 5080 2202 5136 2204
rect 5160 2202 5216 2204
rect 5240 2202 5296 2204
rect 4920 2150 4922 2202
rect 4922 2150 4974 2202
rect 4974 2150 4976 2202
rect 5000 2150 5038 2202
rect 5038 2150 5050 2202
rect 5050 2150 5056 2202
rect 5080 2150 5102 2202
rect 5102 2150 5114 2202
rect 5114 2150 5136 2202
rect 5160 2150 5166 2202
rect 5166 2150 5178 2202
rect 5178 2150 5216 2202
rect 5240 2150 5242 2202
rect 5242 2150 5294 2202
rect 5294 2150 5296 2202
rect 4920 2148 4976 2150
rect 5000 2148 5056 2150
rect 5080 2148 5136 2150
rect 5160 2148 5216 2150
rect 5240 2148 5296 2150
rect 10920 2202 10976 2204
rect 11000 2202 11056 2204
rect 11080 2202 11136 2204
rect 11160 2202 11216 2204
rect 11240 2202 11296 2204
rect 10920 2150 10922 2202
rect 10922 2150 10974 2202
rect 10974 2150 10976 2202
rect 11000 2150 11038 2202
rect 11038 2150 11050 2202
rect 11050 2150 11056 2202
rect 11080 2150 11102 2202
rect 11102 2150 11114 2202
rect 11114 2150 11136 2202
rect 11160 2150 11166 2202
rect 11166 2150 11178 2202
rect 11178 2150 11216 2202
rect 11240 2150 11242 2202
rect 11242 2150 11294 2202
rect 11294 2150 11296 2202
rect 10920 2148 10976 2150
rect 11000 2148 11056 2150
rect 11080 2148 11136 2150
rect 11160 2148 11216 2150
rect 11240 2148 11296 2150
rect 16920 2202 16976 2204
rect 17000 2202 17056 2204
rect 17080 2202 17136 2204
rect 17160 2202 17216 2204
rect 17240 2202 17296 2204
rect 16920 2150 16922 2202
rect 16922 2150 16974 2202
rect 16974 2150 16976 2202
rect 17000 2150 17038 2202
rect 17038 2150 17050 2202
rect 17050 2150 17056 2202
rect 17080 2150 17102 2202
rect 17102 2150 17114 2202
rect 17114 2150 17136 2202
rect 17160 2150 17166 2202
rect 17166 2150 17178 2202
rect 17178 2150 17216 2202
rect 17240 2150 17242 2202
rect 17242 2150 17294 2202
rect 17294 2150 17296 2202
rect 16920 2148 16976 2150
rect 17000 2148 17056 2150
rect 17080 2148 17136 2150
rect 17160 2148 17216 2150
rect 17240 2148 17296 2150
rect 22920 2202 22976 2204
rect 23000 2202 23056 2204
rect 23080 2202 23136 2204
rect 23160 2202 23216 2204
rect 23240 2202 23296 2204
rect 22920 2150 22922 2202
rect 22922 2150 22974 2202
rect 22974 2150 22976 2202
rect 23000 2150 23038 2202
rect 23038 2150 23050 2202
rect 23050 2150 23056 2202
rect 23080 2150 23102 2202
rect 23102 2150 23114 2202
rect 23114 2150 23136 2202
rect 23160 2150 23166 2202
rect 23166 2150 23178 2202
rect 23178 2150 23216 2202
rect 23240 2150 23242 2202
rect 23242 2150 23294 2202
rect 23294 2150 23296 2202
rect 22920 2148 22976 2150
rect 23000 2148 23056 2150
rect 23080 2148 23136 2150
rect 23160 2148 23216 2150
rect 23240 2148 23296 2150
rect 28920 2202 28976 2204
rect 29000 2202 29056 2204
rect 29080 2202 29136 2204
rect 29160 2202 29216 2204
rect 29240 2202 29296 2204
rect 28920 2150 28922 2202
rect 28922 2150 28974 2202
rect 28974 2150 28976 2202
rect 29000 2150 29038 2202
rect 29038 2150 29050 2202
rect 29050 2150 29056 2202
rect 29080 2150 29102 2202
rect 29102 2150 29114 2202
rect 29114 2150 29136 2202
rect 29160 2150 29166 2202
rect 29166 2150 29178 2202
rect 29178 2150 29216 2202
rect 29240 2150 29242 2202
rect 29242 2150 29294 2202
rect 29294 2150 29296 2202
rect 28920 2148 28976 2150
rect 29000 2148 29056 2150
rect 29080 2148 29136 2150
rect 29160 2148 29216 2150
rect 29240 2148 29296 2150
rect 30838 1400 30894 1456
<< metal3 >>
rect 4170 32128 4566 32129
rect 4170 32064 4176 32128
rect 4240 32064 4256 32128
rect 4320 32064 4336 32128
rect 4400 32064 4416 32128
rect 4480 32064 4496 32128
rect 4560 32064 4566 32128
rect 4170 32063 4566 32064
rect 10170 32128 10566 32129
rect 10170 32064 10176 32128
rect 10240 32064 10256 32128
rect 10320 32064 10336 32128
rect 10400 32064 10416 32128
rect 10480 32064 10496 32128
rect 10560 32064 10566 32128
rect 10170 32063 10566 32064
rect 16170 32128 16566 32129
rect 16170 32064 16176 32128
rect 16240 32064 16256 32128
rect 16320 32064 16336 32128
rect 16400 32064 16416 32128
rect 16480 32064 16496 32128
rect 16560 32064 16566 32128
rect 16170 32063 16566 32064
rect 22170 32128 22566 32129
rect 22170 32064 22176 32128
rect 22240 32064 22256 32128
rect 22320 32064 22336 32128
rect 22400 32064 22416 32128
rect 22480 32064 22496 32128
rect 22560 32064 22566 32128
rect 22170 32063 22566 32064
rect 28170 32128 28566 32129
rect 28170 32064 28176 32128
rect 28240 32064 28256 32128
rect 28320 32064 28336 32128
rect 28400 32064 28416 32128
rect 28480 32064 28496 32128
rect 28560 32064 28566 32128
rect 28170 32063 28566 32064
rect 24342 31724 24348 31788
rect 24412 31786 24418 31788
rect 24485 31786 24551 31789
rect 24412 31784 24551 31786
rect 24412 31728 24490 31784
rect 24546 31728 24551 31784
rect 24412 31726 24551 31728
rect 24412 31724 24418 31726
rect 24485 31723 24551 31726
rect 4910 31584 5306 31585
rect 4910 31520 4916 31584
rect 4980 31520 4996 31584
rect 5060 31520 5076 31584
rect 5140 31520 5156 31584
rect 5220 31520 5236 31584
rect 5300 31520 5306 31584
rect 4910 31519 5306 31520
rect 10910 31584 11306 31585
rect 10910 31520 10916 31584
rect 10980 31520 10996 31584
rect 11060 31520 11076 31584
rect 11140 31520 11156 31584
rect 11220 31520 11236 31584
rect 11300 31520 11306 31584
rect 10910 31519 11306 31520
rect 16910 31584 17306 31585
rect 16910 31520 16916 31584
rect 16980 31520 16996 31584
rect 17060 31520 17076 31584
rect 17140 31520 17156 31584
rect 17220 31520 17236 31584
rect 17300 31520 17306 31584
rect 16910 31519 17306 31520
rect 22910 31584 23306 31585
rect 22910 31520 22916 31584
rect 22980 31520 22996 31584
rect 23060 31520 23076 31584
rect 23140 31520 23156 31584
rect 23220 31520 23236 31584
rect 23300 31520 23306 31584
rect 22910 31519 23306 31520
rect 28910 31584 29306 31585
rect 28910 31520 28916 31584
rect 28980 31520 28996 31584
rect 29060 31520 29076 31584
rect 29140 31520 29156 31584
rect 29220 31520 29236 31584
rect 29300 31520 29306 31584
rect 28910 31519 29306 31520
rect 27838 31316 27844 31380
rect 27908 31378 27914 31380
rect 31652 31378 32452 31408
rect 27908 31318 32452 31378
rect 27908 31316 27914 31318
rect 31652 31288 32452 31318
rect 4170 31040 4566 31041
rect 4170 30976 4176 31040
rect 4240 30976 4256 31040
rect 4320 30976 4336 31040
rect 4400 30976 4416 31040
rect 4480 30976 4496 31040
rect 4560 30976 4566 31040
rect 4170 30975 4566 30976
rect 10170 31040 10566 31041
rect 10170 30976 10176 31040
rect 10240 30976 10256 31040
rect 10320 30976 10336 31040
rect 10400 30976 10416 31040
rect 10480 30976 10496 31040
rect 10560 30976 10566 31040
rect 10170 30975 10566 30976
rect 16170 31040 16566 31041
rect 16170 30976 16176 31040
rect 16240 30976 16256 31040
rect 16320 30976 16336 31040
rect 16400 30976 16416 31040
rect 16480 30976 16496 31040
rect 16560 30976 16566 31040
rect 16170 30975 16566 30976
rect 22170 31040 22566 31041
rect 22170 30976 22176 31040
rect 22240 30976 22256 31040
rect 22320 30976 22336 31040
rect 22400 30976 22416 31040
rect 22480 30976 22496 31040
rect 22560 30976 22566 31040
rect 22170 30975 22566 30976
rect 28170 31040 28566 31041
rect 28170 30976 28176 31040
rect 28240 30976 28256 31040
rect 28320 30976 28336 31040
rect 28400 30976 28416 31040
rect 28480 30976 28496 31040
rect 28560 30976 28566 31040
rect 28170 30975 28566 30976
rect 4910 30496 5306 30497
rect 4910 30432 4916 30496
rect 4980 30432 4996 30496
rect 5060 30432 5076 30496
rect 5140 30432 5156 30496
rect 5220 30432 5236 30496
rect 5300 30432 5306 30496
rect 4910 30431 5306 30432
rect 10910 30496 11306 30497
rect 10910 30432 10916 30496
rect 10980 30432 10996 30496
rect 11060 30432 11076 30496
rect 11140 30432 11156 30496
rect 11220 30432 11236 30496
rect 11300 30432 11306 30496
rect 10910 30431 11306 30432
rect 16910 30496 17306 30497
rect 16910 30432 16916 30496
rect 16980 30432 16996 30496
rect 17060 30432 17076 30496
rect 17140 30432 17156 30496
rect 17220 30432 17236 30496
rect 17300 30432 17306 30496
rect 16910 30431 17306 30432
rect 22910 30496 23306 30497
rect 22910 30432 22916 30496
rect 22980 30432 22996 30496
rect 23060 30432 23076 30496
rect 23140 30432 23156 30496
rect 23220 30432 23236 30496
rect 23300 30432 23306 30496
rect 22910 30431 23306 30432
rect 28910 30496 29306 30497
rect 28910 30432 28916 30496
rect 28980 30432 28996 30496
rect 29060 30432 29076 30496
rect 29140 30432 29156 30496
rect 29220 30432 29236 30496
rect 29300 30432 29306 30496
rect 28910 30431 29306 30432
rect 0 30018 800 30048
rect 933 30018 999 30021
rect 0 30016 999 30018
rect 0 29960 938 30016
rect 994 29960 999 30016
rect 0 29958 999 29960
rect 0 29928 800 29958
rect 933 29955 999 29958
rect 4170 29952 4566 29953
rect 4170 29888 4176 29952
rect 4240 29888 4256 29952
rect 4320 29888 4336 29952
rect 4400 29888 4416 29952
rect 4480 29888 4496 29952
rect 4560 29888 4566 29952
rect 4170 29887 4566 29888
rect 10170 29952 10566 29953
rect 10170 29888 10176 29952
rect 10240 29888 10256 29952
rect 10320 29888 10336 29952
rect 10400 29888 10416 29952
rect 10480 29888 10496 29952
rect 10560 29888 10566 29952
rect 10170 29887 10566 29888
rect 16170 29952 16566 29953
rect 16170 29888 16176 29952
rect 16240 29888 16256 29952
rect 16320 29888 16336 29952
rect 16400 29888 16416 29952
rect 16480 29888 16496 29952
rect 16560 29888 16566 29952
rect 16170 29887 16566 29888
rect 22170 29952 22566 29953
rect 22170 29888 22176 29952
rect 22240 29888 22256 29952
rect 22320 29888 22336 29952
rect 22400 29888 22416 29952
rect 22480 29888 22496 29952
rect 22560 29888 22566 29952
rect 22170 29887 22566 29888
rect 28170 29952 28566 29953
rect 28170 29888 28176 29952
rect 28240 29888 28256 29952
rect 28320 29888 28336 29952
rect 28400 29888 28416 29952
rect 28480 29888 28496 29952
rect 28560 29888 28566 29952
rect 28170 29887 28566 29888
rect 4910 29408 5306 29409
rect 4910 29344 4916 29408
rect 4980 29344 4996 29408
rect 5060 29344 5076 29408
rect 5140 29344 5156 29408
rect 5220 29344 5236 29408
rect 5300 29344 5306 29408
rect 4910 29343 5306 29344
rect 10910 29408 11306 29409
rect 10910 29344 10916 29408
rect 10980 29344 10996 29408
rect 11060 29344 11076 29408
rect 11140 29344 11156 29408
rect 11220 29344 11236 29408
rect 11300 29344 11306 29408
rect 10910 29343 11306 29344
rect 16910 29408 17306 29409
rect 16910 29344 16916 29408
rect 16980 29344 16996 29408
rect 17060 29344 17076 29408
rect 17140 29344 17156 29408
rect 17220 29344 17236 29408
rect 17300 29344 17306 29408
rect 16910 29343 17306 29344
rect 22910 29408 23306 29409
rect 22910 29344 22916 29408
rect 22980 29344 22996 29408
rect 23060 29344 23076 29408
rect 23140 29344 23156 29408
rect 23220 29344 23236 29408
rect 23300 29344 23306 29408
rect 22910 29343 23306 29344
rect 28910 29408 29306 29409
rect 28910 29344 28916 29408
rect 28980 29344 28996 29408
rect 29060 29344 29076 29408
rect 29140 29344 29156 29408
rect 29220 29344 29236 29408
rect 29300 29344 29306 29408
rect 28910 29343 29306 29344
rect 4170 28864 4566 28865
rect 4170 28800 4176 28864
rect 4240 28800 4256 28864
rect 4320 28800 4336 28864
rect 4400 28800 4416 28864
rect 4480 28800 4496 28864
rect 4560 28800 4566 28864
rect 4170 28799 4566 28800
rect 10170 28864 10566 28865
rect 10170 28800 10176 28864
rect 10240 28800 10256 28864
rect 10320 28800 10336 28864
rect 10400 28800 10416 28864
rect 10480 28800 10496 28864
rect 10560 28800 10566 28864
rect 10170 28799 10566 28800
rect 16170 28864 16566 28865
rect 16170 28800 16176 28864
rect 16240 28800 16256 28864
rect 16320 28800 16336 28864
rect 16400 28800 16416 28864
rect 16480 28800 16496 28864
rect 16560 28800 16566 28864
rect 16170 28799 16566 28800
rect 22170 28864 22566 28865
rect 22170 28800 22176 28864
rect 22240 28800 22256 28864
rect 22320 28800 22336 28864
rect 22400 28800 22416 28864
rect 22480 28800 22496 28864
rect 22560 28800 22566 28864
rect 22170 28799 22566 28800
rect 28170 28864 28566 28865
rect 28170 28800 28176 28864
rect 28240 28800 28256 28864
rect 28320 28800 28336 28864
rect 28400 28800 28416 28864
rect 28480 28800 28496 28864
rect 28560 28800 28566 28864
rect 28170 28799 28566 28800
rect 4910 28320 5306 28321
rect 4910 28256 4916 28320
rect 4980 28256 4996 28320
rect 5060 28256 5076 28320
rect 5140 28256 5156 28320
rect 5220 28256 5236 28320
rect 5300 28256 5306 28320
rect 4910 28255 5306 28256
rect 10910 28320 11306 28321
rect 10910 28256 10916 28320
rect 10980 28256 10996 28320
rect 11060 28256 11076 28320
rect 11140 28256 11156 28320
rect 11220 28256 11236 28320
rect 11300 28256 11306 28320
rect 10910 28255 11306 28256
rect 16910 28320 17306 28321
rect 16910 28256 16916 28320
rect 16980 28256 16996 28320
rect 17060 28256 17076 28320
rect 17140 28256 17156 28320
rect 17220 28256 17236 28320
rect 17300 28256 17306 28320
rect 16910 28255 17306 28256
rect 22910 28320 23306 28321
rect 22910 28256 22916 28320
rect 22980 28256 22996 28320
rect 23060 28256 23076 28320
rect 23140 28256 23156 28320
rect 23220 28256 23236 28320
rect 23300 28256 23306 28320
rect 22910 28255 23306 28256
rect 28910 28320 29306 28321
rect 28910 28256 28916 28320
rect 28980 28256 28996 28320
rect 29060 28256 29076 28320
rect 29140 28256 29156 28320
rect 29220 28256 29236 28320
rect 29300 28256 29306 28320
rect 28910 28255 29306 28256
rect 22461 27978 22527 27981
rect 23381 27978 23447 27981
rect 22461 27976 23447 27978
rect 22461 27920 22466 27976
rect 22522 27920 23386 27976
rect 23442 27920 23447 27976
rect 22461 27918 23447 27920
rect 22461 27915 22527 27918
rect 23381 27915 23447 27918
rect 4170 27776 4566 27777
rect 4170 27712 4176 27776
rect 4240 27712 4256 27776
rect 4320 27712 4336 27776
rect 4400 27712 4416 27776
rect 4480 27712 4496 27776
rect 4560 27712 4566 27776
rect 4170 27711 4566 27712
rect 10170 27776 10566 27777
rect 10170 27712 10176 27776
rect 10240 27712 10256 27776
rect 10320 27712 10336 27776
rect 10400 27712 10416 27776
rect 10480 27712 10496 27776
rect 10560 27712 10566 27776
rect 10170 27711 10566 27712
rect 16170 27776 16566 27777
rect 16170 27712 16176 27776
rect 16240 27712 16256 27776
rect 16320 27712 16336 27776
rect 16400 27712 16416 27776
rect 16480 27712 16496 27776
rect 16560 27712 16566 27776
rect 16170 27711 16566 27712
rect 22170 27776 22566 27777
rect 22170 27712 22176 27776
rect 22240 27712 22256 27776
rect 22320 27712 22336 27776
rect 22400 27712 22416 27776
rect 22480 27712 22496 27776
rect 22560 27712 22566 27776
rect 22170 27711 22566 27712
rect 28170 27776 28566 27777
rect 28170 27712 28176 27776
rect 28240 27712 28256 27776
rect 28320 27712 28336 27776
rect 28400 27712 28416 27776
rect 28480 27712 28496 27776
rect 28560 27712 28566 27776
rect 28170 27711 28566 27712
rect 24025 27706 24091 27709
rect 24526 27706 24532 27708
rect 24025 27704 24532 27706
rect 24025 27648 24030 27704
rect 24086 27648 24532 27704
rect 24025 27646 24532 27648
rect 24025 27643 24091 27646
rect 24526 27644 24532 27646
rect 24596 27644 24602 27708
rect 4910 27232 5306 27233
rect 4910 27168 4916 27232
rect 4980 27168 4996 27232
rect 5060 27168 5076 27232
rect 5140 27168 5156 27232
rect 5220 27168 5236 27232
rect 5300 27168 5306 27232
rect 4910 27167 5306 27168
rect 10910 27232 11306 27233
rect 10910 27168 10916 27232
rect 10980 27168 10996 27232
rect 11060 27168 11076 27232
rect 11140 27168 11156 27232
rect 11220 27168 11236 27232
rect 11300 27168 11306 27232
rect 10910 27167 11306 27168
rect 16910 27232 17306 27233
rect 16910 27168 16916 27232
rect 16980 27168 16996 27232
rect 17060 27168 17076 27232
rect 17140 27168 17156 27232
rect 17220 27168 17236 27232
rect 17300 27168 17306 27232
rect 16910 27167 17306 27168
rect 22910 27232 23306 27233
rect 22910 27168 22916 27232
rect 22980 27168 22996 27232
rect 23060 27168 23076 27232
rect 23140 27168 23156 27232
rect 23220 27168 23236 27232
rect 23300 27168 23306 27232
rect 22910 27167 23306 27168
rect 28910 27232 29306 27233
rect 28910 27168 28916 27232
rect 28980 27168 28996 27232
rect 29060 27168 29076 27232
rect 29140 27168 29156 27232
rect 29220 27168 29236 27232
rect 29300 27168 29306 27232
rect 28910 27167 29306 27168
rect 4170 26688 4566 26689
rect 4170 26624 4176 26688
rect 4240 26624 4256 26688
rect 4320 26624 4336 26688
rect 4400 26624 4416 26688
rect 4480 26624 4496 26688
rect 4560 26624 4566 26688
rect 4170 26623 4566 26624
rect 10170 26688 10566 26689
rect 10170 26624 10176 26688
rect 10240 26624 10256 26688
rect 10320 26624 10336 26688
rect 10400 26624 10416 26688
rect 10480 26624 10496 26688
rect 10560 26624 10566 26688
rect 10170 26623 10566 26624
rect 16170 26688 16566 26689
rect 16170 26624 16176 26688
rect 16240 26624 16256 26688
rect 16320 26624 16336 26688
rect 16400 26624 16416 26688
rect 16480 26624 16496 26688
rect 16560 26624 16566 26688
rect 16170 26623 16566 26624
rect 22170 26688 22566 26689
rect 22170 26624 22176 26688
rect 22240 26624 22256 26688
rect 22320 26624 22336 26688
rect 22400 26624 22416 26688
rect 22480 26624 22496 26688
rect 22560 26624 22566 26688
rect 22170 26623 22566 26624
rect 28170 26688 28566 26689
rect 28170 26624 28176 26688
rect 28240 26624 28256 26688
rect 28320 26624 28336 26688
rect 28400 26624 28416 26688
rect 28480 26624 28496 26688
rect 28560 26624 28566 26688
rect 28170 26623 28566 26624
rect 18689 26348 18755 26349
rect 18638 26284 18644 26348
rect 18708 26346 18755 26348
rect 18708 26344 18800 26346
rect 18750 26288 18800 26344
rect 18708 26286 18800 26288
rect 18708 26284 18755 26286
rect 18689 26283 18755 26284
rect 4910 26144 5306 26145
rect 4910 26080 4916 26144
rect 4980 26080 4996 26144
rect 5060 26080 5076 26144
rect 5140 26080 5156 26144
rect 5220 26080 5236 26144
rect 5300 26080 5306 26144
rect 4910 26079 5306 26080
rect 10910 26144 11306 26145
rect 10910 26080 10916 26144
rect 10980 26080 10996 26144
rect 11060 26080 11076 26144
rect 11140 26080 11156 26144
rect 11220 26080 11236 26144
rect 11300 26080 11306 26144
rect 10910 26079 11306 26080
rect 16910 26144 17306 26145
rect 16910 26080 16916 26144
rect 16980 26080 16996 26144
rect 17060 26080 17076 26144
rect 17140 26080 17156 26144
rect 17220 26080 17236 26144
rect 17300 26080 17306 26144
rect 16910 26079 17306 26080
rect 22910 26144 23306 26145
rect 22910 26080 22916 26144
rect 22980 26080 22996 26144
rect 23060 26080 23076 26144
rect 23140 26080 23156 26144
rect 23220 26080 23236 26144
rect 23300 26080 23306 26144
rect 22910 26079 23306 26080
rect 28910 26144 29306 26145
rect 28910 26080 28916 26144
rect 28980 26080 28996 26144
rect 29060 26080 29076 26144
rect 29140 26080 29156 26144
rect 29220 26080 29236 26144
rect 29300 26080 29306 26144
rect 28910 26079 29306 26080
rect 4170 25600 4566 25601
rect 4170 25536 4176 25600
rect 4240 25536 4256 25600
rect 4320 25536 4336 25600
rect 4400 25536 4416 25600
rect 4480 25536 4496 25600
rect 4560 25536 4566 25600
rect 4170 25535 4566 25536
rect 10170 25600 10566 25601
rect 10170 25536 10176 25600
rect 10240 25536 10256 25600
rect 10320 25536 10336 25600
rect 10400 25536 10416 25600
rect 10480 25536 10496 25600
rect 10560 25536 10566 25600
rect 10170 25535 10566 25536
rect 16170 25600 16566 25601
rect 16170 25536 16176 25600
rect 16240 25536 16256 25600
rect 16320 25536 16336 25600
rect 16400 25536 16416 25600
rect 16480 25536 16496 25600
rect 16560 25536 16566 25600
rect 16170 25535 16566 25536
rect 22170 25600 22566 25601
rect 22170 25536 22176 25600
rect 22240 25536 22256 25600
rect 22320 25536 22336 25600
rect 22400 25536 22416 25600
rect 22480 25536 22496 25600
rect 22560 25536 22566 25600
rect 22170 25535 22566 25536
rect 28170 25600 28566 25601
rect 28170 25536 28176 25600
rect 28240 25536 28256 25600
rect 28320 25536 28336 25600
rect 28400 25536 28416 25600
rect 28480 25536 28496 25600
rect 28560 25536 28566 25600
rect 28170 25535 28566 25536
rect 31293 25258 31359 25261
rect 31652 25258 32452 25288
rect 31293 25256 32452 25258
rect 31293 25200 31298 25256
rect 31354 25200 32452 25256
rect 31293 25198 32452 25200
rect 31293 25195 31359 25198
rect 31652 25168 32452 25198
rect 4910 25056 5306 25057
rect 4910 24992 4916 25056
rect 4980 24992 4996 25056
rect 5060 24992 5076 25056
rect 5140 24992 5156 25056
rect 5220 24992 5236 25056
rect 5300 24992 5306 25056
rect 4910 24991 5306 24992
rect 10910 25056 11306 25057
rect 10910 24992 10916 25056
rect 10980 24992 10996 25056
rect 11060 24992 11076 25056
rect 11140 24992 11156 25056
rect 11220 24992 11236 25056
rect 11300 24992 11306 25056
rect 10910 24991 11306 24992
rect 16910 25056 17306 25057
rect 16910 24992 16916 25056
rect 16980 24992 16996 25056
rect 17060 24992 17076 25056
rect 17140 24992 17156 25056
rect 17220 24992 17236 25056
rect 17300 24992 17306 25056
rect 16910 24991 17306 24992
rect 22910 25056 23306 25057
rect 22910 24992 22916 25056
rect 22980 24992 22996 25056
rect 23060 24992 23076 25056
rect 23140 24992 23156 25056
rect 23220 24992 23236 25056
rect 23300 24992 23306 25056
rect 22910 24991 23306 24992
rect 28910 25056 29306 25057
rect 28910 24992 28916 25056
rect 28980 24992 28996 25056
rect 29060 24992 29076 25056
rect 29140 24992 29156 25056
rect 29220 24992 29236 25056
rect 29300 24992 29306 25056
rect 28910 24991 29306 24992
rect 4170 24512 4566 24513
rect 4170 24448 4176 24512
rect 4240 24448 4256 24512
rect 4320 24448 4336 24512
rect 4400 24448 4416 24512
rect 4480 24448 4496 24512
rect 4560 24448 4566 24512
rect 4170 24447 4566 24448
rect 10170 24512 10566 24513
rect 10170 24448 10176 24512
rect 10240 24448 10256 24512
rect 10320 24448 10336 24512
rect 10400 24448 10416 24512
rect 10480 24448 10496 24512
rect 10560 24448 10566 24512
rect 10170 24447 10566 24448
rect 16170 24512 16566 24513
rect 16170 24448 16176 24512
rect 16240 24448 16256 24512
rect 16320 24448 16336 24512
rect 16400 24448 16416 24512
rect 16480 24448 16496 24512
rect 16560 24448 16566 24512
rect 16170 24447 16566 24448
rect 22170 24512 22566 24513
rect 22170 24448 22176 24512
rect 22240 24448 22256 24512
rect 22320 24448 22336 24512
rect 22400 24448 22416 24512
rect 22480 24448 22496 24512
rect 22560 24448 22566 24512
rect 22170 24447 22566 24448
rect 28170 24512 28566 24513
rect 28170 24448 28176 24512
rect 28240 24448 28256 24512
rect 28320 24448 28336 24512
rect 28400 24448 28416 24512
rect 28480 24448 28496 24512
rect 28560 24448 28566 24512
rect 28170 24447 28566 24448
rect 4910 23968 5306 23969
rect 0 23898 800 23928
rect 4910 23904 4916 23968
rect 4980 23904 4996 23968
rect 5060 23904 5076 23968
rect 5140 23904 5156 23968
rect 5220 23904 5236 23968
rect 5300 23904 5306 23968
rect 4910 23903 5306 23904
rect 10910 23968 11306 23969
rect 10910 23904 10916 23968
rect 10980 23904 10996 23968
rect 11060 23904 11076 23968
rect 11140 23904 11156 23968
rect 11220 23904 11236 23968
rect 11300 23904 11306 23968
rect 10910 23903 11306 23904
rect 16910 23968 17306 23969
rect 16910 23904 16916 23968
rect 16980 23904 16996 23968
rect 17060 23904 17076 23968
rect 17140 23904 17156 23968
rect 17220 23904 17236 23968
rect 17300 23904 17306 23968
rect 16910 23903 17306 23904
rect 22910 23968 23306 23969
rect 22910 23904 22916 23968
rect 22980 23904 22996 23968
rect 23060 23904 23076 23968
rect 23140 23904 23156 23968
rect 23220 23904 23236 23968
rect 23300 23904 23306 23968
rect 22910 23903 23306 23904
rect 28910 23968 29306 23969
rect 28910 23904 28916 23968
rect 28980 23904 28996 23968
rect 29060 23904 29076 23968
rect 29140 23904 29156 23968
rect 29220 23904 29236 23968
rect 29300 23904 29306 23968
rect 28910 23903 29306 23904
rect 933 23898 999 23901
rect 0 23896 999 23898
rect 0 23840 938 23896
rect 994 23840 999 23896
rect 0 23838 999 23840
rect 0 23808 800 23838
rect 933 23835 999 23838
rect 10685 23626 10751 23629
rect 15326 23626 15332 23628
rect 10685 23624 15332 23626
rect 10685 23568 10690 23624
rect 10746 23568 15332 23624
rect 10685 23566 15332 23568
rect 10685 23563 10751 23566
rect 15326 23564 15332 23566
rect 15396 23626 15402 23628
rect 17217 23626 17283 23629
rect 15396 23624 17283 23626
rect 15396 23568 17222 23624
rect 17278 23568 17283 23624
rect 15396 23566 17283 23568
rect 15396 23564 15402 23566
rect 17217 23563 17283 23566
rect 17861 23490 17927 23493
rect 19333 23490 19399 23493
rect 17861 23488 19399 23490
rect 17861 23432 17866 23488
rect 17922 23432 19338 23488
rect 19394 23432 19399 23488
rect 17861 23430 19399 23432
rect 17861 23427 17927 23430
rect 19333 23427 19399 23430
rect 4170 23424 4566 23425
rect 4170 23360 4176 23424
rect 4240 23360 4256 23424
rect 4320 23360 4336 23424
rect 4400 23360 4416 23424
rect 4480 23360 4496 23424
rect 4560 23360 4566 23424
rect 4170 23359 4566 23360
rect 10170 23424 10566 23425
rect 10170 23360 10176 23424
rect 10240 23360 10256 23424
rect 10320 23360 10336 23424
rect 10400 23360 10416 23424
rect 10480 23360 10496 23424
rect 10560 23360 10566 23424
rect 10170 23359 10566 23360
rect 16170 23424 16566 23425
rect 16170 23360 16176 23424
rect 16240 23360 16256 23424
rect 16320 23360 16336 23424
rect 16400 23360 16416 23424
rect 16480 23360 16496 23424
rect 16560 23360 16566 23424
rect 16170 23359 16566 23360
rect 22170 23424 22566 23425
rect 22170 23360 22176 23424
rect 22240 23360 22256 23424
rect 22320 23360 22336 23424
rect 22400 23360 22416 23424
rect 22480 23360 22496 23424
rect 22560 23360 22566 23424
rect 22170 23359 22566 23360
rect 28170 23424 28566 23425
rect 28170 23360 28176 23424
rect 28240 23360 28256 23424
rect 28320 23360 28336 23424
rect 28400 23360 28416 23424
rect 28480 23360 28496 23424
rect 28560 23360 28566 23424
rect 28170 23359 28566 23360
rect 10225 23082 10291 23085
rect 12617 23082 12683 23085
rect 10225 23080 12683 23082
rect 10225 23024 10230 23080
rect 10286 23024 12622 23080
rect 12678 23024 12683 23080
rect 10225 23022 12683 23024
rect 10225 23019 10291 23022
rect 12617 23019 12683 23022
rect 4910 22880 5306 22881
rect 4910 22816 4916 22880
rect 4980 22816 4996 22880
rect 5060 22816 5076 22880
rect 5140 22816 5156 22880
rect 5220 22816 5236 22880
rect 5300 22816 5306 22880
rect 4910 22815 5306 22816
rect 10910 22880 11306 22881
rect 10910 22816 10916 22880
rect 10980 22816 10996 22880
rect 11060 22816 11076 22880
rect 11140 22816 11156 22880
rect 11220 22816 11236 22880
rect 11300 22816 11306 22880
rect 10910 22815 11306 22816
rect 16910 22880 17306 22881
rect 16910 22816 16916 22880
rect 16980 22816 16996 22880
rect 17060 22816 17076 22880
rect 17140 22816 17156 22880
rect 17220 22816 17236 22880
rect 17300 22816 17306 22880
rect 16910 22815 17306 22816
rect 22910 22880 23306 22881
rect 22910 22816 22916 22880
rect 22980 22816 22996 22880
rect 23060 22816 23076 22880
rect 23140 22816 23156 22880
rect 23220 22816 23236 22880
rect 23300 22816 23306 22880
rect 22910 22815 23306 22816
rect 28910 22880 29306 22881
rect 28910 22816 28916 22880
rect 28980 22816 28996 22880
rect 29060 22816 29076 22880
rect 29140 22816 29156 22880
rect 29220 22816 29236 22880
rect 29300 22816 29306 22880
rect 28910 22815 29306 22816
rect 4170 22336 4566 22337
rect 4170 22272 4176 22336
rect 4240 22272 4256 22336
rect 4320 22272 4336 22336
rect 4400 22272 4416 22336
rect 4480 22272 4496 22336
rect 4560 22272 4566 22336
rect 4170 22271 4566 22272
rect 10170 22336 10566 22337
rect 10170 22272 10176 22336
rect 10240 22272 10256 22336
rect 10320 22272 10336 22336
rect 10400 22272 10416 22336
rect 10480 22272 10496 22336
rect 10560 22272 10566 22336
rect 10170 22271 10566 22272
rect 16170 22336 16566 22337
rect 16170 22272 16176 22336
rect 16240 22272 16256 22336
rect 16320 22272 16336 22336
rect 16400 22272 16416 22336
rect 16480 22272 16496 22336
rect 16560 22272 16566 22336
rect 16170 22271 16566 22272
rect 22170 22336 22566 22337
rect 22170 22272 22176 22336
rect 22240 22272 22256 22336
rect 22320 22272 22336 22336
rect 22400 22272 22416 22336
rect 22480 22272 22496 22336
rect 22560 22272 22566 22336
rect 22170 22271 22566 22272
rect 28170 22336 28566 22337
rect 28170 22272 28176 22336
rect 28240 22272 28256 22336
rect 28320 22272 28336 22336
rect 28400 22272 28416 22336
rect 28480 22272 28496 22336
rect 28560 22272 28566 22336
rect 28170 22271 28566 22272
rect 16481 21994 16547 21997
rect 17401 21994 17467 21997
rect 16481 21992 17467 21994
rect 16481 21936 16486 21992
rect 16542 21936 17406 21992
rect 17462 21936 17467 21992
rect 16481 21934 17467 21936
rect 16481 21931 16547 21934
rect 17401 21931 17467 21934
rect 20989 21994 21055 21997
rect 24342 21994 24348 21996
rect 20989 21992 24348 21994
rect 20989 21936 20994 21992
rect 21050 21936 24348 21992
rect 20989 21934 24348 21936
rect 20989 21931 21055 21934
rect 24342 21932 24348 21934
rect 24412 21932 24418 21996
rect 4910 21792 5306 21793
rect 4910 21728 4916 21792
rect 4980 21728 4996 21792
rect 5060 21728 5076 21792
rect 5140 21728 5156 21792
rect 5220 21728 5236 21792
rect 5300 21728 5306 21792
rect 4910 21727 5306 21728
rect 10910 21792 11306 21793
rect 10910 21728 10916 21792
rect 10980 21728 10996 21792
rect 11060 21728 11076 21792
rect 11140 21728 11156 21792
rect 11220 21728 11236 21792
rect 11300 21728 11306 21792
rect 10910 21727 11306 21728
rect 16910 21792 17306 21793
rect 16910 21728 16916 21792
rect 16980 21728 16996 21792
rect 17060 21728 17076 21792
rect 17140 21728 17156 21792
rect 17220 21728 17236 21792
rect 17300 21728 17306 21792
rect 16910 21727 17306 21728
rect 22910 21792 23306 21793
rect 22910 21728 22916 21792
rect 22980 21728 22996 21792
rect 23060 21728 23076 21792
rect 23140 21728 23156 21792
rect 23220 21728 23236 21792
rect 23300 21728 23306 21792
rect 22910 21727 23306 21728
rect 28910 21792 29306 21793
rect 28910 21728 28916 21792
rect 28980 21728 28996 21792
rect 29060 21728 29076 21792
rect 29140 21728 29156 21792
rect 29220 21728 29236 21792
rect 29300 21728 29306 21792
rect 28910 21727 29306 21728
rect 4170 21248 4566 21249
rect 4170 21184 4176 21248
rect 4240 21184 4256 21248
rect 4320 21184 4336 21248
rect 4400 21184 4416 21248
rect 4480 21184 4496 21248
rect 4560 21184 4566 21248
rect 4170 21183 4566 21184
rect 10170 21248 10566 21249
rect 10170 21184 10176 21248
rect 10240 21184 10256 21248
rect 10320 21184 10336 21248
rect 10400 21184 10416 21248
rect 10480 21184 10496 21248
rect 10560 21184 10566 21248
rect 10170 21183 10566 21184
rect 16170 21248 16566 21249
rect 16170 21184 16176 21248
rect 16240 21184 16256 21248
rect 16320 21184 16336 21248
rect 16400 21184 16416 21248
rect 16480 21184 16496 21248
rect 16560 21184 16566 21248
rect 16170 21183 16566 21184
rect 22170 21248 22566 21249
rect 22170 21184 22176 21248
rect 22240 21184 22256 21248
rect 22320 21184 22336 21248
rect 22400 21184 22416 21248
rect 22480 21184 22496 21248
rect 22560 21184 22566 21248
rect 22170 21183 22566 21184
rect 28170 21248 28566 21249
rect 28170 21184 28176 21248
rect 28240 21184 28256 21248
rect 28320 21184 28336 21248
rect 28400 21184 28416 21248
rect 28480 21184 28496 21248
rect 28560 21184 28566 21248
rect 28170 21183 28566 21184
rect 9673 21042 9739 21045
rect 10317 21042 10383 21045
rect 19333 21042 19399 21045
rect 9673 21040 19399 21042
rect 9673 20984 9678 21040
rect 9734 20984 10322 21040
rect 10378 20984 19338 21040
rect 19394 20984 19399 21040
rect 9673 20982 19399 20984
rect 9673 20979 9739 20982
rect 10317 20979 10383 20982
rect 19333 20979 19399 20982
rect 10593 20906 10659 20909
rect 16941 20906 17007 20909
rect 10593 20904 17007 20906
rect 10593 20848 10598 20904
rect 10654 20848 16946 20904
rect 17002 20848 17007 20904
rect 10593 20846 17007 20848
rect 10593 20843 10659 20846
rect 16941 20843 17007 20846
rect 4910 20704 5306 20705
rect 4910 20640 4916 20704
rect 4980 20640 4996 20704
rect 5060 20640 5076 20704
rect 5140 20640 5156 20704
rect 5220 20640 5236 20704
rect 5300 20640 5306 20704
rect 4910 20639 5306 20640
rect 10910 20704 11306 20705
rect 10910 20640 10916 20704
rect 10980 20640 10996 20704
rect 11060 20640 11076 20704
rect 11140 20640 11156 20704
rect 11220 20640 11236 20704
rect 11300 20640 11306 20704
rect 10910 20639 11306 20640
rect 16910 20704 17306 20705
rect 16910 20640 16916 20704
rect 16980 20640 16996 20704
rect 17060 20640 17076 20704
rect 17140 20640 17156 20704
rect 17220 20640 17236 20704
rect 17300 20640 17306 20704
rect 16910 20639 17306 20640
rect 22910 20704 23306 20705
rect 22910 20640 22916 20704
rect 22980 20640 22996 20704
rect 23060 20640 23076 20704
rect 23140 20640 23156 20704
rect 23220 20640 23236 20704
rect 23300 20640 23306 20704
rect 22910 20639 23306 20640
rect 28910 20704 29306 20705
rect 28910 20640 28916 20704
rect 28980 20640 28996 20704
rect 29060 20640 29076 20704
rect 29140 20640 29156 20704
rect 29220 20640 29236 20704
rect 29300 20640 29306 20704
rect 28910 20639 29306 20640
rect 4170 20160 4566 20161
rect 4170 20096 4176 20160
rect 4240 20096 4256 20160
rect 4320 20096 4336 20160
rect 4400 20096 4416 20160
rect 4480 20096 4496 20160
rect 4560 20096 4566 20160
rect 4170 20095 4566 20096
rect 10170 20160 10566 20161
rect 10170 20096 10176 20160
rect 10240 20096 10256 20160
rect 10320 20096 10336 20160
rect 10400 20096 10416 20160
rect 10480 20096 10496 20160
rect 10560 20096 10566 20160
rect 10170 20095 10566 20096
rect 16170 20160 16566 20161
rect 16170 20096 16176 20160
rect 16240 20096 16256 20160
rect 16320 20096 16336 20160
rect 16400 20096 16416 20160
rect 16480 20096 16496 20160
rect 16560 20096 16566 20160
rect 16170 20095 16566 20096
rect 22170 20160 22566 20161
rect 22170 20096 22176 20160
rect 22240 20096 22256 20160
rect 22320 20096 22336 20160
rect 22400 20096 22416 20160
rect 22480 20096 22496 20160
rect 22560 20096 22566 20160
rect 22170 20095 22566 20096
rect 28170 20160 28566 20161
rect 28170 20096 28176 20160
rect 28240 20096 28256 20160
rect 28320 20096 28336 20160
rect 28400 20096 28416 20160
rect 28480 20096 28496 20160
rect 28560 20096 28566 20160
rect 28170 20095 28566 20096
rect 15929 19954 15995 19957
rect 20069 19954 20135 19957
rect 24485 19954 24551 19957
rect 15929 19952 16130 19954
rect 15929 19896 15934 19952
rect 15990 19896 16130 19952
rect 15929 19894 16130 19896
rect 15929 19891 15995 19894
rect 4910 19616 5306 19617
rect 4910 19552 4916 19616
rect 4980 19552 4996 19616
rect 5060 19552 5076 19616
rect 5140 19552 5156 19616
rect 5220 19552 5236 19616
rect 5300 19552 5306 19616
rect 4910 19551 5306 19552
rect 10910 19616 11306 19617
rect 10910 19552 10916 19616
rect 10980 19552 10996 19616
rect 11060 19552 11076 19616
rect 11140 19552 11156 19616
rect 11220 19552 11236 19616
rect 11300 19552 11306 19616
rect 10910 19551 11306 19552
rect 15469 19410 15535 19413
rect 16070 19410 16130 19894
rect 20069 19952 24551 19954
rect 20069 19896 20074 19952
rect 20130 19896 24490 19952
rect 24546 19896 24551 19952
rect 20069 19894 24551 19896
rect 20069 19891 20135 19894
rect 24485 19891 24551 19894
rect 19333 19818 19399 19821
rect 19885 19818 19951 19821
rect 19333 19816 19951 19818
rect 19333 19760 19338 19816
rect 19394 19760 19890 19816
rect 19946 19760 19951 19816
rect 19333 19758 19951 19760
rect 19333 19755 19399 19758
rect 19885 19755 19951 19758
rect 16910 19616 17306 19617
rect 16910 19552 16916 19616
rect 16980 19552 16996 19616
rect 17060 19552 17076 19616
rect 17140 19552 17156 19616
rect 17220 19552 17236 19616
rect 17300 19552 17306 19616
rect 16910 19551 17306 19552
rect 22910 19616 23306 19617
rect 22910 19552 22916 19616
rect 22980 19552 22996 19616
rect 23060 19552 23076 19616
rect 23140 19552 23156 19616
rect 23220 19552 23236 19616
rect 23300 19552 23306 19616
rect 22910 19551 23306 19552
rect 28910 19616 29306 19617
rect 28910 19552 28916 19616
rect 28980 19552 28996 19616
rect 29060 19552 29076 19616
rect 29140 19552 29156 19616
rect 29220 19552 29236 19616
rect 29300 19552 29306 19616
rect 28910 19551 29306 19552
rect 16941 19410 17007 19413
rect 20621 19410 20687 19413
rect 15469 19408 20687 19410
rect 15469 19352 15474 19408
rect 15530 19352 16946 19408
rect 17002 19352 20626 19408
rect 20682 19352 20687 19408
rect 15469 19350 20687 19352
rect 15469 19347 15535 19350
rect 16941 19347 17007 19350
rect 20621 19347 20687 19350
rect 30925 19138 30991 19141
rect 31652 19138 32452 19168
rect 30925 19136 32452 19138
rect 30925 19080 30930 19136
rect 30986 19080 32452 19136
rect 30925 19078 32452 19080
rect 30925 19075 30991 19078
rect 4170 19072 4566 19073
rect 4170 19008 4176 19072
rect 4240 19008 4256 19072
rect 4320 19008 4336 19072
rect 4400 19008 4416 19072
rect 4480 19008 4496 19072
rect 4560 19008 4566 19072
rect 4170 19007 4566 19008
rect 10170 19072 10566 19073
rect 10170 19008 10176 19072
rect 10240 19008 10256 19072
rect 10320 19008 10336 19072
rect 10400 19008 10416 19072
rect 10480 19008 10496 19072
rect 10560 19008 10566 19072
rect 10170 19007 10566 19008
rect 16170 19072 16566 19073
rect 16170 19008 16176 19072
rect 16240 19008 16256 19072
rect 16320 19008 16336 19072
rect 16400 19008 16416 19072
rect 16480 19008 16496 19072
rect 16560 19008 16566 19072
rect 16170 19007 16566 19008
rect 22170 19072 22566 19073
rect 22170 19008 22176 19072
rect 22240 19008 22256 19072
rect 22320 19008 22336 19072
rect 22400 19008 22416 19072
rect 22480 19008 22496 19072
rect 22560 19008 22566 19072
rect 22170 19007 22566 19008
rect 28170 19072 28566 19073
rect 28170 19008 28176 19072
rect 28240 19008 28256 19072
rect 28320 19008 28336 19072
rect 28400 19008 28416 19072
rect 28480 19008 28496 19072
rect 28560 19008 28566 19072
rect 31652 19048 32452 19078
rect 28170 19007 28566 19008
rect 16297 18866 16363 18869
rect 18229 18866 18295 18869
rect 16297 18864 18295 18866
rect 16297 18808 16302 18864
rect 16358 18808 18234 18864
rect 18290 18808 18295 18864
rect 16297 18806 18295 18808
rect 16297 18803 16363 18806
rect 18229 18803 18295 18806
rect 14733 18730 14799 18733
rect 17953 18730 18019 18733
rect 14733 18728 18019 18730
rect 14733 18672 14738 18728
rect 14794 18672 17958 18728
rect 18014 18672 18019 18728
rect 14733 18670 18019 18672
rect 14733 18667 14799 18670
rect 17953 18667 18019 18670
rect 4910 18528 5306 18529
rect 4910 18464 4916 18528
rect 4980 18464 4996 18528
rect 5060 18464 5076 18528
rect 5140 18464 5156 18528
rect 5220 18464 5236 18528
rect 5300 18464 5306 18528
rect 4910 18463 5306 18464
rect 10910 18528 11306 18529
rect 10910 18464 10916 18528
rect 10980 18464 10996 18528
rect 11060 18464 11076 18528
rect 11140 18464 11156 18528
rect 11220 18464 11236 18528
rect 11300 18464 11306 18528
rect 10910 18463 11306 18464
rect 16910 18528 17306 18529
rect 16910 18464 16916 18528
rect 16980 18464 16996 18528
rect 17060 18464 17076 18528
rect 17140 18464 17156 18528
rect 17220 18464 17236 18528
rect 17300 18464 17306 18528
rect 16910 18463 17306 18464
rect 22910 18528 23306 18529
rect 22910 18464 22916 18528
rect 22980 18464 22996 18528
rect 23060 18464 23076 18528
rect 23140 18464 23156 18528
rect 23220 18464 23236 18528
rect 23300 18464 23306 18528
rect 22910 18463 23306 18464
rect 28910 18528 29306 18529
rect 28910 18464 28916 18528
rect 28980 18464 28996 18528
rect 29060 18464 29076 18528
rect 29140 18464 29156 18528
rect 29220 18464 29236 18528
rect 29300 18464 29306 18528
rect 28910 18463 29306 18464
rect 4170 17984 4566 17985
rect 4170 17920 4176 17984
rect 4240 17920 4256 17984
rect 4320 17920 4336 17984
rect 4400 17920 4416 17984
rect 4480 17920 4496 17984
rect 4560 17920 4566 17984
rect 4170 17919 4566 17920
rect 10170 17984 10566 17985
rect 10170 17920 10176 17984
rect 10240 17920 10256 17984
rect 10320 17920 10336 17984
rect 10400 17920 10416 17984
rect 10480 17920 10496 17984
rect 10560 17920 10566 17984
rect 10170 17919 10566 17920
rect 16170 17984 16566 17985
rect 16170 17920 16176 17984
rect 16240 17920 16256 17984
rect 16320 17920 16336 17984
rect 16400 17920 16416 17984
rect 16480 17920 16496 17984
rect 16560 17920 16566 17984
rect 16170 17919 16566 17920
rect 22170 17984 22566 17985
rect 22170 17920 22176 17984
rect 22240 17920 22256 17984
rect 22320 17920 22336 17984
rect 22400 17920 22416 17984
rect 22480 17920 22496 17984
rect 22560 17920 22566 17984
rect 22170 17919 22566 17920
rect 28170 17984 28566 17985
rect 28170 17920 28176 17984
rect 28240 17920 28256 17984
rect 28320 17920 28336 17984
rect 28400 17920 28416 17984
rect 28480 17920 28496 17984
rect 28560 17920 28566 17984
rect 28170 17919 28566 17920
rect 1393 17914 1459 17917
rect 798 17912 1459 17914
rect 798 17856 1398 17912
rect 1454 17856 1459 17912
rect 798 17854 1459 17856
rect 798 17808 858 17854
rect 1393 17851 1459 17854
rect 0 17718 858 17808
rect 12249 17778 12315 17781
rect 15193 17778 15259 17781
rect 12249 17776 15259 17778
rect 12249 17720 12254 17776
rect 12310 17720 15198 17776
rect 15254 17720 15259 17776
rect 12249 17718 15259 17720
rect 0 17688 800 17718
rect 12249 17715 12315 17718
rect 15193 17715 15259 17718
rect 15929 17778 15995 17781
rect 18689 17778 18755 17781
rect 15929 17776 18755 17778
rect 15929 17720 15934 17776
rect 15990 17720 18694 17776
rect 18750 17720 18755 17776
rect 15929 17718 18755 17720
rect 15929 17715 15995 17718
rect 18689 17715 18755 17718
rect 9581 17642 9647 17645
rect 15653 17642 15719 17645
rect 17309 17642 17375 17645
rect 9581 17640 17375 17642
rect 9581 17584 9586 17640
rect 9642 17584 15658 17640
rect 15714 17584 17314 17640
rect 17370 17584 17375 17640
rect 9581 17582 17375 17584
rect 9581 17579 9647 17582
rect 15653 17579 15719 17582
rect 17309 17579 17375 17582
rect 19333 17642 19399 17645
rect 21081 17642 21147 17645
rect 19333 17640 21147 17642
rect 19333 17584 19338 17640
rect 19394 17584 21086 17640
rect 21142 17584 21147 17640
rect 19333 17582 21147 17584
rect 19333 17579 19399 17582
rect 21081 17579 21147 17582
rect 4910 17440 5306 17441
rect 4910 17376 4916 17440
rect 4980 17376 4996 17440
rect 5060 17376 5076 17440
rect 5140 17376 5156 17440
rect 5220 17376 5236 17440
rect 5300 17376 5306 17440
rect 4910 17375 5306 17376
rect 10910 17440 11306 17441
rect 10910 17376 10916 17440
rect 10980 17376 10996 17440
rect 11060 17376 11076 17440
rect 11140 17376 11156 17440
rect 11220 17376 11236 17440
rect 11300 17376 11306 17440
rect 10910 17375 11306 17376
rect 16910 17440 17306 17441
rect 16910 17376 16916 17440
rect 16980 17376 16996 17440
rect 17060 17376 17076 17440
rect 17140 17376 17156 17440
rect 17220 17376 17236 17440
rect 17300 17376 17306 17440
rect 16910 17375 17306 17376
rect 22910 17440 23306 17441
rect 22910 17376 22916 17440
rect 22980 17376 22996 17440
rect 23060 17376 23076 17440
rect 23140 17376 23156 17440
rect 23220 17376 23236 17440
rect 23300 17376 23306 17440
rect 22910 17375 23306 17376
rect 28910 17440 29306 17441
rect 28910 17376 28916 17440
rect 28980 17376 28996 17440
rect 29060 17376 29076 17440
rect 29140 17376 29156 17440
rect 29220 17376 29236 17440
rect 29300 17376 29306 17440
rect 28910 17375 29306 17376
rect 11421 17370 11487 17373
rect 14457 17370 14523 17373
rect 11421 17368 14523 17370
rect 11421 17312 11426 17368
rect 11482 17312 14462 17368
rect 14518 17312 14523 17368
rect 11421 17310 14523 17312
rect 11421 17307 11487 17310
rect 14457 17307 14523 17310
rect 15193 17370 15259 17373
rect 15326 17370 15332 17372
rect 15193 17368 15332 17370
rect 15193 17312 15198 17368
rect 15254 17312 15332 17368
rect 15193 17310 15332 17312
rect 15193 17307 15259 17310
rect 15326 17308 15332 17310
rect 15396 17308 15402 17372
rect 10869 17234 10935 17237
rect 14733 17234 14799 17237
rect 10869 17232 14799 17234
rect 10869 17176 10874 17232
rect 10930 17176 14738 17232
rect 14794 17176 14799 17232
rect 10869 17174 14799 17176
rect 10869 17171 10935 17174
rect 14733 17171 14799 17174
rect 16481 17234 16547 17237
rect 27838 17234 27844 17236
rect 16481 17232 27844 17234
rect 16481 17176 16486 17232
rect 16542 17176 27844 17232
rect 16481 17174 27844 17176
rect 16481 17171 16547 17174
rect 27838 17172 27844 17174
rect 27908 17172 27914 17236
rect 8017 17098 8083 17101
rect 13445 17098 13511 17101
rect 8017 17096 13511 17098
rect 8017 17040 8022 17096
rect 8078 17040 13450 17096
rect 13506 17040 13511 17096
rect 8017 17038 13511 17040
rect 8017 17035 8083 17038
rect 13445 17035 13511 17038
rect 4170 16896 4566 16897
rect 4170 16832 4176 16896
rect 4240 16832 4256 16896
rect 4320 16832 4336 16896
rect 4400 16832 4416 16896
rect 4480 16832 4496 16896
rect 4560 16832 4566 16896
rect 4170 16831 4566 16832
rect 10170 16896 10566 16897
rect 10170 16832 10176 16896
rect 10240 16832 10256 16896
rect 10320 16832 10336 16896
rect 10400 16832 10416 16896
rect 10480 16832 10496 16896
rect 10560 16832 10566 16896
rect 10170 16831 10566 16832
rect 16170 16896 16566 16897
rect 16170 16832 16176 16896
rect 16240 16832 16256 16896
rect 16320 16832 16336 16896
rect 16400 16832 16416 16896
rect 16480 16832 16496 16896
rect 16560 16832 16566 16896
rect 16170 16831 16566 16832
rect 22170 16896 22566 16897
rect 22170 16832 22176 16896
rect 22240 16832 22256 16896
rect 22320 16832 22336 16896
rect 22400 16832 22416 16896
rect 22480 16832 22496 16896
rect 22560 16832 22566 16896
rect 22170 16831 22566 16832
rect 28170 16896 28566 16897
rect 28170 16832 28176 16896
rect 28240 16832 28256 16896
rect 28320 16832 28336 16896
rect 28400 16832 28416 16896
rect 28480 16832 28496 16896
rect 28560 16832 28566 16896
rect 28170 16831 28566 16832
rect 4910 16352 5306 16353
rect 4910 16288 4916 16352
rect 4980 16288 4996 16352
rect 5060 16288 5076 16352
rect 5140 16288 5156 16352
rect 5220 16288 5236 16352
rect 5300 16288 5306 16352
rect 4910 16287 5306 16288
rect 10910 16352 11306 16353
rect 10910 16288 10916 16352
rect 10980 16288 10996 16352
rect 11060 16288 11076 16352
rect 11140 16288 11156 16352
rect 11220 16288 11236 16352
rect 11300 16288 11306 16352
rect 10910 16287 11306 16288
rect 16910 16352 17306 16353
rect 16910 16288 16916 16352
rect 16980 16288 16996 16352
rect 17060 16288 17076 16352
rect 17140 16288 17156 16352
rect 17220 16288 17236 16352
rect 17300 16288 17306 16352
rect 16910 16287 17306 16288
rect 22910 16352 23306 16353
rect 22910 16288 22916 16352
rect 22980 16288 22996 16352
rect 23060 16288 23076 16352
rect 23140 16288 23156 16352
rect 23220 16288 23236 16352
rect 23300 16288 23306 16352
rect 22910 16287 23306 16288
rect 28910 16352 29306 16353
rect 28910 16288 28916 16352
rect 28980 16288 28996 16352
rect 29060 16288 29076 16352
rect 29140 16288 29156 16352
rect 29220 16288 29236 16352
rect 29300 16288 29306 16352
rect 28910 16287 29306 16288
rect 19609 16282 19675 16285
rect 20989 16282 21055 16285
rect 19609 16280 21055 16282
rect 19609 16224 19614 16280
rect 19670 16224 20994 16280
rect 21050 16224 21055 16280
rect 19609 16222 21055 16224
rect 19609 16219 19675 16222
rect 20989 16219 21055 16222
rect 4170 15808 4566 15809
rect 4170 15744 4176 15808
rect 4240 15744 4256 15808
rect 4320 15744 4336 15808
rect 4400 15744 4416 15808
rect 4480 15744 4496 15808
rect 4560 15744 4566 15808
rect 4170 15743 4566 15744
rect 10170 15808 10566 15809
rect 10170 15744 10176 15808
rect 10240 15744 10256 15808
rect 10320 15744 10336 15808
rect 10400 15744 10416 15808
rect 10480 15744 10496 15808
rect 10560 15744 10566 15808
rect 10170 15743 10566 15744
rect 16170 15808 16566 15809
rect 16170 15744 16176 15808
rect 16240 15744 16256 15808
rect 16320 15744 16336 15808
rect 16400 15744 16416 15808
rect 16480 15744 16496 15808
rect 16560 15744 16566 15808
rect 16170 15743 16566 15744
rect 22170 15808 22566 15809
rect 22170 15744 22176 15808
rect 22240 15744 22256 15808
rect 22320 15744 22336 15808
rect 22400 15744 22416 15808
rect 22480 15744 22496 15808
rect 22560 15744 22566 15808
rect 22170 15743 22566 15744
rect 28170 15808 28566 15809
rect 28170 15744 28176 15808
rect 28240 15744 28256 15808
rect 28320 15744 28336 15808
rect 28400 15744 28416 15808
rect 28480 15744 28496 15808
rect 28560 15744 28566 15808
rect 28170 15743 28566 15744
rect 4910 15264 5306 15265
rect 4910 15200 4916 15264
rect 4980 15200 4996 15264
rect 5060 15200 5076 15264
rect 5140 15200 5156 15264
rect 5220 15200 5236 15264
rect 5300 15200 5306 15264
rect 4910 15199 5306 15200
rect 10910 15264 11306 15265
rect 10910 15200 10916 15264
rect 10980 15200 10996 15264
rect 11060 15200 11076 15264
rect 11140 15200 11156 15264
rect 11220 15200 11236 15264
rect 11300 15200 11306 15264
rect 10910 15199 11306 15200
rect 16910 15264 17306 15265
rect 16910 15200 16916 15264
rect 16980 15200 16996 15264
rect 17060 15200 17076 15264
rect 17140 15200 17156 15264
rect 17220 15200 17236 15264
rect 17300 15200 17306 15264
rect 16910 15199 17306 15200
rect 22910 15264 23306 15265
rect 22910 15200 22916 15264
rect 22980 15200 22996 15264
rect 23060 15200 23076 15264
rect 23140 15200 23156 15264
rect 23220 15200 23236 15264
rect 23300 15200 23306 15264
rect 22910 15199 23306 15200
rect 28910 15264 29306 15265
rect 28910 15200 28916 15264
rect 28980 15200 28996 15264
rect 29060 15200 29076 15264
rect 29140 15200 29156 15264
rect 29220 15200 29236 15264
rect 29300 15200 29306 15264
rect 28910 15199 29306 15200
rect 24393 15194 24459 15197
rect 24526 15194 24532 15196
rect 24393 15192 24532 15194
rect 24393 15136 24398 15192
rect 24454 15136 24532 15192
rect 24393 15134 24532 15136
rect 24393 15131 24459 15134
rect 24526 15132 24532 15134
rect 24596 15132 24602 15196
rect 4170 14720 4566 14721
rect 4170 14656 4176 14720
rect 4240 14656 4256 14720
rect 4320 14656 4336 14720
rect 4400 14656 4416 14720
rect 4480 14656 4496 14720
rect 4560 14656 4566 14720
rect 4170 14655 4566 14656
rect 10170 14720 10566 14721
rect 10170 14656 10176 14720
rect 10240 14656 10256 14720
rect 10320 14656 10336 14720
rect 10400 14656 10416 14720
rect 10480 14656 10496 14720
rect 10560 14656 10566 14720
rect 10170 14655 10566 14656
rect 16170 14720 16566 14721
rect 16170 14656 16176 14720
rect 16240 14656 16256 14720
rect 16320 14656 16336 14720
rect 16400 14656 16416 14720
rect 16480 14656 16496 14720
rect 16560 14656 16566 14720
rect 16170 14655 16566 14656
rect 22170 14720 22566 14721
rect 22170 14656 22176 14720
rect 22240 14656 22256 14720
rect 22320 14656 22336 14720
rect 22400 14656 22416 14720
rect 22480 14656 22496 14720
rect 22560 14656 22566 14720
rect 22170 14655 22566 14656
rect 28170 14720 28566 14721
rect 28170 14656 28176 14720
rect 28240 14656 28256 14720
rect 28320 14656 28336 14720
rect 28400 14656 28416 14720
rect 28480 14656 28496 14720
rect 28560 14656 28566 14720
rect 28170 14655 28566 14656
rect 4910 14176 5306 14177
rect 4910 14112 4916 14176
rect 4980 14112 4996 14176
rect 5060 14112 5076 14176
rect 5140 14112 5156 14176
rect 5220 14112 5236 14176
rect 5300 14112 5306 14176
rect 4910 14111 5306 14112
rect 10910 14176 11306 14177
rect 10910 14112 10916 14176
rect 10980 14112 10996 14176
rect 11060 14112 11076 14176
rect 11140 14112 11156 14176
rect 11220 14112 11236 14176
rect 11300 14112 11306 14176
rect 10910 14111 11306 14112
rect 16910 14176 17306 14177
rect 16910 14112 16916 14176
rect 16980 14112 16996 14176
rect 17060 14112 17076 14176
rect 17140 14112 17156 14176
rect 17220 14112 17236 14176
rect 17300 14112 17306 14176
rect 16910 14111 17306 14112
rect 22910 14176 23306 14177
rect 22910 14112 22916 14176
rect 22980 14112 22996 14176
rect 23060 14112 23076 14176
rect 23140 14112 23156 14176
rect 23220 14112 23236 14176
rect 23300 14112 23306 14176
rect 22910 14111 23306 14112
rect 28910 14176 29306 14177
rect 28910 14112 28916 14176
rect 28980 14112 28996 14176
rect 29060 14112 29076 14176
rect 29140 14112 29156 14176
rect 29220 14112 29236 14176
rect 29300 14112 29306 14176
rect 28910 14111 29306 14112
rect 4170 13632 4566 13633
rect 4170 13568 4176 13632
rect 4240 13568 4256 13632
rect 4320 13568 4336 13632
rect 4400 13568 4416 13632
rect 4480 13568 4496 13632
rect 4560 13568 4566 13632
rect 4170 13567 4566 13568
rect 10170 13632 10566 13633
rect 10170 13568 10176 13632
rect 10240 13568 10256 13632
rect 10320 13568 10336 13632
rect 10400 13568 10416 13632
rect 10480 13568 10496 13632
rect 10560 13568 10566 13632
rect 10170 13567 10566 13568
rect 16170 13632 16566 13633
rect 16170 13568 16176 13632
rect 16240 13568 16256 13632
rect 16320 13568 16336 13632
rect 16400 13568 16416 13632
rect 16480 13568 16496 13632
rect 16560 13568 16566 13632
rect 16170 13567 16566 13568
rect 22170 13632 22566 13633
rect 22170 13568 22176 13632
rect 22240 13568 22256 13632
rect 22320 13568 22336 13632
rect 22400 13568 22416 13632
rect 22480 13568 22496 13632
rect 22560 13568 22566 13632
rect 22170 13567 22566 13568
rect 28170 13632 28566 13633
rect 28170 13568 28176 13632
rect 28240 13568 28256 13632
rect 28320 13568 28336 13632
rect 28400 13568 28416 13632
rect 28480 13568 28496 13632
rect 28560 13568 28566 13632
rect 28170 13567 28566 13568
rect 4910 13088 5306 13089
rect 4910 13024 4916 13088
rect 4980 13024 4996 13088
rect 5060 13024 5076 13088
rect 5140 13024 5156 13088
rect 5220 13024 5236 13088
rect 5300 13024 5306 13088
rect 4910 13023 5306 13024
rect 10910 13088 11306 13089
rect 10910 13024 10916 13088
rect 10980 13024 10996 13088
rect 11060 13024 11076 13088
rect 11140 13024 11156 13088
rect 11220 13024 11236 13088
rect 11300 13024 11306 13088
rect 10910 13023 11306 13024
rect 16910 13088 17306 13089
rect 16910 13024 16916 13088
rect 16980 13024 16996 13088
rect 17060 13024 17076 13088
rect 17140 13024 17156 13088
rect 17220 13024 17236 13088
rect 17300 13024 17306 13088
rect 16910 13023 17306 13024
rect 22910 13088 23306 13089
rect 22910 13024 22916 13088
rect 22980 13024 22996 13088
rect 23060 13024 23076 13088
rect 23140 13024 23156 13088
rect 23220 13024 23236 13088
rect 23300 13024 23306 13088
rect 22910 13023 23306 13024
rect 28910 13088 29306 13089
rect 28910 13024 28916 13088
rect 28980 13024 28996 13088
rect 29060 13024 29076 13088
rect 29140 13024 29156 13088
rect 29220 13024 29236 13088
rect 29300 13024 29306 13088
rect 28910 13023 29306 13024
rect 31293 13018 31359 13021
rect 31652 13018 32452 13048
rect 31293 13016 32452 13018
rect 31293 12960 31298 13016
rect 31354 12960 32452 13016
rect 31293 12958 32452 12960
rect 31293 12955 31359 12958
rect 31652 12928 32452 12958
rect 10501 12882 10567 12885
rect 15326 12882 15332 12884
rect 10501 12880 15332 12882
rect 10501 12824 10506 12880
rect 10562 12824 15332 12880
rect 10501 12822 15332 12824
rect 10501 12819 10567 12822
rect 15326 12820 15332 12822
rect 15396 12820 15402 12884
rect 4170 12544 4566 12545
rect 4170 12480 4176 12544
rect 4240 12480 4256 12544
rect 4320 12480 4336 12544
rect 4400 12480 4416 12544
rect 4480 12480 4496 12544
rect 4560 12480 4566 12544
rect 4170 12479 4566 12480
rect 10170 12544 10566 12545
rect 10170 12480 10176 12544
rect 10240 12480 10256 12544
rect 10320 12480 10336 12544
rect 10400 12480 10416 12544
rect 10480 12480 10496 12544
rect 10560 12480 10566 12544
rect 10170 12479 10566 12480
rect 16170 12544 16566 12545
rect 16170 12480 16176 12544
rect 16240 12480 16256 12544
rect 16320 12480 16336 12544
rect 16400 12480 16416 12544
rect 16480 12480 16496 12544
rect 16560 12480 16566 12544
rect 16170 12479 16566 12480
rect 22170 12544 22566 12545
rect 22170 12480 22176 12544
rect 22240 12480 22256 12544
rect 22320 12480 22336 12544
rect 22400 12480 22416 12544
rect 22480 12480 22496 12544
rect 22560 12480 22566 12544
rect 22170 12479 22566 12480
rect 28170 12544 28566 12545
rect 28170 12480 28176 12544
rect 28240 12480 28256 12544
rect 28320 12480 28336 12544
rect 28400 12480 28416 12544
rect 28480 12480 28496 12544
rect 28560 12480 28566 12544
rect 28170 12479 28566 12480
rect 23197 12202 23263 12205
rect 23197 12200 23490 12202
rect 23197 12144 23202 12200
rect 23258 12144 23490 12200
rect 23197 12142 23490 12144
rect 23197 12139 23263 12142
rect 4910 12000 5306 12001
rect 4910 11936 4916 12000
rect 4980 11936 4996 12000
rect 5060 11936 5076 12000
rect 5140 11936 5156 12000
rect 5220 11936 5236 12000
rect 5300 11936 5306 12000
rect 4910 11935 5306 11936
rect 10910 12000 11306 12001
rect 10910 11936 10916 12000
rect 10980 11936 10996 12000
rect 11060 11936 11076 12000
rect 11140 11936 11156 12000
rect 11220 11936 11236 12000
rect 11300 11936 11306 12000
rect 10910 11935 11306 11936
rect 16910 12000 17306 12001
rect 16910 11936 16916 12000
rect 16980 11936 16996 12000
rect 17060 11936 17076 12000
rect 17140 11936 17156 12000
rect 17220 11936 17236 12000
rect 17300 11936 17306 12000
rect 16910 11935 17306 11936
rect 22910 12000 23306 12001
rect 22910 11936 22916 12000
rect 22980 11936 22996 12000
rect 23060 11936 23076 12000
rect 23140 11936 23156 12000
rect 23220 11936 23236 12000
rect 23300 11936 23306 12000
rect 22910 11935 23306 11936
rect 23430 11930 23490 12142
rect 28910 12000 29306 12001
rect 28910 11936 28916 12000
rect 28980 11936 28996 12000
rect 29060 11936 29076 12000
rect 29140 11936 29156 12000
rect 29220 11936 29236 12000
rect 29300 11936 29306 12000
rect 28910 11935 29306 11936
rect 23565 11930 23631 11933
rect 23430 11928 23631 11930
rect 23430 11872 23570 11928
rect 23626 11872 23631 11928
rect 23430 11870 23631 11872
rect 23565 11867 23631 11870
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4170 11456 4566 11457
rect 4170 11392 4176 11456
rect 4240 11392 4256 11456
rect 4320 11392 4336 11456
rect 4400 11392 4416 11456
rect 4480 11392 4496 11456
rect 4560 11392 4566 11456
rect 4170 11391 4566 11392
rect 10170 11456 10566 11457
rect 10170 11392 10176 11456
rect 10240 11392 10256 11456
rect 10320 11392 10336 11456
rect 10400 11392 10416 11456
rect 10480 11392 10496 11456
rect 10560 11392 10566 11456
rect 10170 11391 10566 11392
rect 16170 11456 16566 11457
rect 16170 11392 16176 11456
rect 16240 11392 16256 11456
rect 16320 11392 16336 11456
rect 16400 11392 16416 11456
rect 16480 11392 16496 11456
rect 16560 11392 16566 11456
rect 16170 11391 16566 11392
rect 22170 11456 22566 11457
rect 22170 11392 22176 11456
rect 22240 11392 22256 11456
rect 22320 11392 22336 11456
rect 22400 11392 22416 11456
rect 22480 11392 22496 11456
rect 22560 11392 22566 11456
rect 22170 11391 22566 11392
rect 28170 11456 28566 11457
rect 28170 11392 28176 11456
rect 28240 11392 28256 11456
rect 28320 11392 28336 11456
rect 28400 11392 28416 11456
rect 28480 11392 28496 11456
rect 28560 11392 28566 11456
rect 28170 11391 28566 11392
rect 15377 11116 15443 11117
rect 15326 11114 15332 11116
rect 15286 11054 15332 11114
rect 15396 11112 15443 11116
rect 15438 11056 15443 11112
rect 15326 11052 15332 11054
rect 15396 11052 15443 11056
rect 15377 11051 15443 11052
rect 4910 10912 5306 10913
rect 4910 10848 4916 10912
rect 4980 10848 4996 10912
rect 5060 10848 5076 10912
rect 5140 10848 5156 10912
rect 5220 10848 5236 10912
rect 5300 10848 5306 10912
rect 4910 10847 5306 10848
rect 10910 10912 11306 10913
rect 10910 10848 10916 10912
rect 10980 10848 10996 10912
rect 11060 10848 11076 10912
rect 11140 10848 11156 10912
rect 11220 10848 11236 10912
rect 11300 10848 11306 10912
rect 10910 10847 11306 10848
rect 16910 10912 17306 10913
rect 16910 10848 16916 10912
rect 16980 10848 16996 10912
rect 17060 10848 17076 10912
rect 17140 10848 17156 10912
rect 17220 10848 17236 10912
rect 17300 10848 17306 10912
rect 16910 10847 17306 10848
rect 22910 10912 23306 10913
rect 22910 10848 22916 10912
rect 22980 10848 22996 10912
rect 23060 10848 23076 10912
rect 23140 10848 23156 10912
rect 23220 10848 23236 10912
rect 23300 10848 23306 10912
rect 22910 10847 23306 10848
rect 28910 10912 29306 10913
rect 28910 10848 28916 10912
rect 28980 10848 28996 10912
rect 29060 10848 29076 10912
rect 29140 10848 29156 10912
rect 29220 10848 29236 10912
rect 29300 10848 29306 10912
rect 28910 10847 29306 10848
rect 4170 10368 4566 10369
rect 4170 10304 4176 10368
rect 4240 10304 4256 10368
rect 4320 10304 4336 10368
rect 4400 10304 4416 10368
rect 4480 10304 4496 10368
rect 4560 10304 4566 10368
rect 4170 10303 4566 10304
rect 10170 10368 10566 10369
rect 10170 10304 10176 10368
rect 10240 10304 10256 10368
rect 10320 10304 10336 10368
rect 10400 10304 10416 10368
rect 10480 10304 10496 10368
rect 10560 10304 10566 10368
rect 10170 10303 10566 10304
rect 16170 10368 16566 10369
rect 16170 10304 16176 10368
rect 16240 10304 16256 10368
rect 16320 10304 16336 10368
rect 16400 10304 16416 10368
rect 16480 10304 16496 10368
rect 16560 10304 16566 10368
rect 16170 10303 16566 10304
rect 22170 10368 22566 10369
rect 22170 10304 22176 10368
rect 22240 10304 22256 10368
rect 22320 10304 22336 10368
rect 22400 10304 22416 10368
rect 22480 10304 22496 10368
rect 22560 10304 22566 10368
rect 22170 10303 22566 10304
rect 28170 10368 28566 10369
rect 28170 10304 28176 10368
rect 28240 10304 28256 10368
rect 28320 10304 28336 10368
rect 28400 10304 28416 10368
rect 28480 10304 28496 10368
rect 28560 10304 28566 10368
rect 28170 10303 28566 10304
rect 23013 10026 23079 10029
rect 23013 10024 23490 10026
rect 23013 9968 23018 10024
rect 23074 9968 23490 10024
rect 23013 9966 23490 9968
rect 23013 9963 23079 9966
rect 4910 9824 5306 9825
rect 4910 9760 4916 9824
rect 4980 9760 4996 9824
rect 5060 9760 5076 9824
rect 5140 9760 5156 9824
rect 5220 9760 5236 9824
rect 5300 9760 5306 9824
rect 4910 9759 5306 9760
rect 10910 9824 11306 9825
rect 10910 9760 10916 9824
rect 10980 9760 10996 9824
rect 11060 9760 11076 9824
rect 11140 9760 11156 9824
rect 11220 9760 11236 9824
rect 11300 9760 11306 9824
rect 10910 9759 11306 9760
rect 16910 9824 17306 9825
rect 16910 9760 16916 9824
rect 16980 9760 16996 9824
rect 17060 9760 17076 9824
rect 17140 9760 17156 9824
rect 17220 9760 17236 9824
rect 17300 9760 17306 9824
rect 16910 9759 17306 9760
rect 22910 9824 23306 9825
rect 22910 9760 22916 9824
rect 22980 9760 22996 9824
rect 23060 9760 23076 9824
rect 23140 9760 23156 9824
rect 23220 9760 23236 9824
rect 23300 9760 23306 9824
rect 22910 9759 23306 9760
rect 22553 9754 22619 9757
rect 22553 9752 22754 9754
rect 22553 9696 22558 9752
rect 22614 9696 22754 9752
rect 22553 9694 22754 9696
rect 22553 9691 22619 9694
rect 22694 9693 22754 9694
rect 22694 9688 22803 9693
rect 22694 9632 22742 9688
rect 22798 9632 22803 9688
rect 22694 9630 22803 9632
rect 22737 9627 22803 9630
rect 23289 9690 23355 9693
rect 23430 9690 23490 9966
rect 28910 9824 29306 9825
rect 28910 9760 28916 9824
rect 28980 9760 28996 9824
rect 29060 9760 29076 9824
rect 29140 9760 29156 9824
rect 29220 9760 29236 9824
rect 29300 9760 29306 9824
rect 28910 9759 29306 9760
rect 23289 9688 23490 9690
rect 23289 9632 23294 9688
rect 23350 9632 23490 9688
rect 23289 9630 23490 9632
rect 23289 9627 23355 9630
rect 4170 9280 4566 9281
rect 4170 9216 4176 9280
rect 4240 9216 4256 9280
rect 4320 9216 4336 9280
rect 4400 9216 4416 9280
rect 4480 9216 4496 9280
rect 4560 9216 4566 9280
rect 4170 9215 4566 9216
rect 10170 9280 10566 9281
rect 10170 9216 10176 9280
rect 10240 9216 10256 9280
rect 10320 9216 10336 9280
rect 10400 9216 10416 9280
rect 10480 9216 10496 9280
rect 10560 9216 10566 9280
rect 10170 9215 10566 9216
rect 16170 9280 16566 9281
rect 16170 9216 16176 9280
rect 16240 9216 16256 9280
rect 16320 9216 16336 9280
rect 16400 9216 16416 9280
rect 16480 9216 16496 9280
rect 16560 9216 16566 9280
rect 16170 9215 16566 9216
rect 22170 9280 22566 9281
rect 22170 9216 22176 9280
rect 22240 9216 22256 9280
rect 22320 9216 22336 9280
rect 22400 9216 22416 9280
rect 22480 9216 22496 9280
rect 22560 9216 22566 9280
rect 22170 9215 22566 9216
rect 28170 9280 28566 9281
rect 28170 9216 28176 9280
rect 28240 9216 28256 9280
rect 28320 9216 28336 9280
rect 28400 9216 28416 9280
rect 28480 9216 28496 9280
rect 28560 9216 28566 9280
rect 28170 9215 28566 9216
rect 23289 8938 23355 8941
rect 25129 8938 25195 8941
rect 23289 8936 25195 8938
rect 23289 8880 23294 8936
rect 23350 8880 25134 8936
rect 25190 8880 25195 8936
rect 23289 8878 25195 8880
rect 23289 8875 23355 8878
rect 25129 8875 25195 8878
rect 17861 8802 17927 8805
rect 18638 8802 18644 8804
rect 17861 8800 18644 8802
rect 17861 8744 17866 8800
rect 17922 8744 18644 8800
rect 17861 8742 18644 8744
rect 17861 8739 17927 8742
rect 18638 8740 18644 8742
rect 18708 8740 18714 8804
rect 4910 8736 5306 8737
rect 4910 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5306 8736
rect 4910 8671 5306 8672
rect 10910 8736 11306 8737
rect 10910 8672 10916 8736
rect 10980 8672 10996 8736
rect 11060 8672 11076 8736
rect 11140 8672 11156 8736
rect 11220 8672 11236 8736
rect 11300 8672 11306 8736
rect 10910 8671 11306 8672
rect 16910 8736 17306 8737
rect 16910 8672 16916 8736
rect 16980 8672 16996 8736
rect 17060 8672 17076 8736
rect 17140 8672 17156 8736
rect 17220 8672 17236 8736
rect 17300 8672 17306 8736
rect 16910 8671 17306 8672
rect 22910 8736 23306 8737
rect 22910 8672 22916 8736
rect 22980 8672 22996 8736
rect 23060 8672 23076 8736
rect 23140 8672 23156 8736
rect 23220 8672 23236 8736
rect 23300 8672 23306 8736
rect 22910 8671 23306 8672
rect 28910 8736 29306 8737
rect 28910 8672 28916 8736
rect 28980 8672 28996 8736
rect 29060 8672 29076 8736
rect 29140 8672 29156 8736
rect 29220 8672 29236 8736
rect 29300 8672 29306 8736
rect 28910 8671 29306 8672
rect 4170 8192 4566 8193
rect 4170 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4566 8192
rect 4170 8127 4566 8128
rect 10170 8192 10566 8193
rect 10170 8128 10176 8192
rect 10240 8128 10256 8192
rect 10320 8128 10336 8192
rect 10400 8128 10416 8192
rect 10480 8128 10496 8192
rect 10560 8128 10566 8192
rect 10170 8127 10566 8128
rect 16170 8192 16566 8193
rect 16170 8128 16176 8192
rect 16240 8128 16256 8192
rect 16320 8128 16336 8192
rect 16400 8128 16416 8192
rect 16480 8128 16496 8192
rect 16560 8128 16566 8192
rect 16170 8127 16566 8128
rect 22170 8192 22566 8193
rect 22170 8128 22176 8192
rect 22240 8128 22256 8192
rect 22320 8128 22336 8192
rect 22400 8128 22416 8192
rect 22480 8128 22496 8192
rect 22560 8128 22566 8192
rect 22170 8127 22566 8128
rect 28170 8192 28566 8193
rect 28170 8128 28176 8192
rect 28240 8128 28256 8192
rect 28320 8128 28336 8192
rect 28400 8128 28416 8192
rect 28480 8128 28496 8192
rect 28560 8128 28566 8192
rect 28170 8127 28566 8128
rect 4910 7648 5306 7649
rect 4910 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5306 7648
rect 4910 7583 5306 7584
rect 10910 7648 11306 7649
rect 10910 7584 10916 7648
rect 10980 7584 10996 7648
rect 11060 7584 11076 7648
rect 11140 7584 11156 7648
rect 11220 7584 11236 7648
rect 11300 7584 11306 7648
rect 10910 7583 11306 7584
rect 16910 7648 17306 7649
rect 16910 7584 16916 7648
rect 16980 7584 16996 7648
rect 17060 7584 17076 7648
rect 17140 7584 17156 7648
rect 17220 7584 17236 7648
rect 17300 7584 17306 7648
rect 16910 7583 17306 7584
rect 22910 7648 23306 7649
rect 22910 7584 22916 7648
rect 22980 7584 22996 7648
rect 23060 7584 23076 7648
rect 23140 7584 23156 7648
rect 23220 7584 23236 7648
rect 23300 7584 23306 7648
rect 22910 7583 23306 7584
rect 28910 7648 29306 7649
rect 28910 7584 28916 7648
rect 28980 7584 28996 7648
rect 29060 7584 29076 7648
rect 29140 7584 29156 7648
rect 29220 7584 29236 7648
rect 29300 7584 29306 7648
rect 28910 7583 29306 7584
rect 31293 7578 31359 7581
rect 31652 7578 32452 7608
rect 31293 7576 32452 7578
rect 31293 7520 31298 7576
rect 31354 7520 32452 7576
rect 31293 7518 32452 7520
rect 31293 7515 31359 7518
rect 31652 7488 32452 7518
rect 4170 7104 4566 7105
rect 4170 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4566 7104
rect 4170 7039 4566 7040
rect 10170 7104 10566 7105
rect 10170 7040 10176 7104
rect 10240 7040 10256 7104
rect 10320 7040 10336 7104
rect 10400 7040 10416 7104
rect 10480 7040 10496 7104
rect 10560 7040 10566 7104
rect 10170 7039 10566 7040
rect 16170 7104 16566 7105
rect 16170 7040 16176 7104
rect 16240 7040 16256 7104
rect 16320 7040 16336 7104
rect 16400 7040 16416 7104
rect 16480 7040 16496 7104
rect 16560 7040 16566 7104
rect 16170 7039 16566 7040
rect 22170 7104 22566 7105
rect 22170 7040 22176 7104
rect 22240 7040 22256 7104
rect 22320 7040 22336 7104
rect 22400 7040 22416 7104
rect 22480 7040 22496 7104
rect 22560 7040 22566 7104
rect 22170 7039 22566 7040
rect 28170 7104 28566 7105
rect 28170 7040 28176 7104
rect 28240 7040 28256 7104
rect 28320 7040 28336 7104
rect 28400 7040 28416 7104
rect 28480 7040 28496 7104
rect 28560 7040 28566 7104
rect 28170 7039 28566 7040
rect 4910 6560 5306 6561
rect 4910 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5306 6560
rect 4910 6495 5306 6496
rect 10910 6560 11306 6561
rect 10910 6496 10916 6560
rect 10980 6496 10996 6560
rect 11060 6496 11076 6560
rect 11140 6496 11156 6560
rect 11220 6496 11236 6560
rect 11300 6496 11306 6560
rect 10910 6495 11306 6496
rect 16910 6560 17306 6561
rect 16910 6496 16916 6560
rect 16980 6496 16996 6560
rect 17060 6496 17076 6560
rect 17140 6496 17156 6560
rect 17220 6496 17236 6560
rect 17300 6496 17306 6560
rect 16910 6495 17306 6496
rect 22910 6560 23306 6561
rect 22910 6496 22916 6560
rect 22980 6496 22996 6560
rect 23060 6496 23076 6560
rect 23140 6496 23156 6560
rect 23220 6496 23236 6560
rect 23300 6496 23306 6560
rect 22910 6495 23306 6496
rect 28910 6560 29306 6561
rect 28910 6496 28916 6560
rect 28980 6496 28996 6560
rect 29060 6496 29076 6560
rect 29140 6496 29156 6560
rect 29220 6496 29236 6560
rect 29300 6496 29306 6560
rect 28910 6495 29306 6496
rect 4170 6016 4566 6017
rect 4170 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4566 6016
rect 4170 5951 4566 5952
rect 10170 6016 10566 6017
rect 10170 5952 10176 6016
rect 10240 5952 10256 6016
rect 10320 5952 10336 6016
rect 10400 5952 10416 6016
rect 10480 5952 10496 6016
rect 10560 5952 10566 6016
rect 10170 5951 10566 5952
rect 16170 6016 16566 6017
rect 16170 5952 16176 6016
rect 16240 5952 16256 6016
rect 16320 5952 16336 6016
rect 16400 5952 16416 6016
rect 16480 5952 16496 6016
rect 16560 5952 16566 6016
rect 16170 5951 16566 5952
rect 22170 6016 22566 6017
rect 22170 5952 22176 6016
rect 22240 5952 22256 6016
rect 22320 5952 22336 6016
rect 22400 5952 22416 6016
rect 22480 5952 22496 6016
rect 22560 5952 22566 6016
rect 22170 5951 22566 5952
rect 28170 6016 28566 6017
rect 28170 5952 28176 6016
rect 28240 5952 28256 6016
rect 28320 5952 28336 6016
rect 28400 5952 28416 6016
rect 28480 5952 28496 6016
rect 28560 5952 28566 6016
rect 28170 5951 28566 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 4910 5472 5306 5473
rect 4910 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5306 5472
rect 4910 5407 5306 5408
rect 10910 5472 11306 5473
rect 10910 5408 10916 5472
rect 10980 5408 10996 5472
rect 11060 5408 11076 5472
rect 11140 5408 11156 5472
rect 11220 5408 11236 5472
rect 11300 5408 11306 5472
rect 10910 5407 11306 5408
rect 16910 5472 17306 5473
rect 16910 5408 16916 5472
rect 16980 5408 16996 5472
rect 17060 5408 17076 5472
rect 17140 5408 17156 5472
rect 17220 5408 17236 5472
rect 17300 5408 17306 5472
rect 16910 5407 17306 5408
rect 22910 5472 23306 5473
rect 22910 5408 22916 5472
rect 22980 5408 22996 5472
rect 23060 5408 23076 5472
rect 23140 5408 23156 5472
rect 23220 5408 23236 5472
rect 23300 5408 23306 5472
rect 22910 5407 23306 5408
rect 28910 5472 29306 5473
rect 28910 5408 28916 5472
rect 28980 5408 28996 5472
rect 29060 5408 29076 5472
rect 29140 5408 29156 5472
rect 29220 5408 29236 5472
rect 29300 5408 29306 5472
rect 28910 5407 29306 5408
rect 4170 4928 4566 4929
rect 4170 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4566 4928
rect 4170 4863 4566 4864
rect 10170 4928 10566 4929
rect 10170 4864 10176 4928
rect 10240 4864 10256 4928
rect 10320 4864 10336 4928
rect 10400 4864 10416 4928
rect 10480 4864 10496 4928
rect 10560 4864 10566 4928
rect 10170 4863 10566 4864
rect 16170 4928 16566 4929
rect 16170 4864 16176 4928
rect 16240 4864 16256 4928
rect 16320 4864 16336 4928
rect 16400 4864 16416 4928
rect 16480 4864 16496 4928
rect 16560 4864 16566 4928
rect 16170 4863 16566 4864
rect 22170 4928 22566 4929
rect 22170 4864 22176 4928
rect 22240 4864 22256 4928
rect 22320 4864 22336 4928
rect 22400 4864 22416 4928
rect 22480 4864 22496 4928
rect 22560 4864 22566 4928
rect 22170 4863 22566 4864
rect 28170 4928 28566 4929
rect 28170 4864 28176 4928
rect 28240 4864 28256 4928
rect 28320 4864 28336 4928
rect 28400 4864 28416 4928
rect 28480 4864 28496 4928
rect 28560 4864 28566 4928
rect 28170 4863 28566 4864
rect 4910 4384 5306 4385
rect 4910 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5306 4384
rect 4910 4319 5306 4320
rect 10910 4384 11306 4385
rect 10910 4320 10916 4384
rect 10980 4320 10996 4384
rect 11060 4320 11076 4384
rect 11140 4320 11156 4384
rect 11220 4320 11236 4384
rect 11300 4320 11306 4384
rect 10910 4319 11306 4320
rect 16910 4384 17306 4385
rect 16910 4320 16916 4384
rect 16980 4320 16996 4384
rect 17060 4320 17076 4384
rect 17140 4320 17156 4384
rect 17220 4320 17236 4384
rect 17300 4320 17306 4384
rect 16910 4319 17306 4320
rect 22910 4384 23306 4385
rect 22910 4320 22916 4384
rect 22980 4320 22996 4384
rect 23060 4320 23076 4384
rect 23140 4320 23156 4384
rect 23220 4320 23236 4384
rect 23300 4320 23306 4384
rect 22910 4319 23306 4320
rect 28910 4384 29306 4385
rect 28910 4320 28916 4384
rect 28980 4320 28996 4384
rect 29060 4320 29076 4384
rect 29140 4320 29156 4384
rect 29220 4320 29236 4384
rect 29300 4320 29306 4384
rect 28910 4319 29306 4320
rect 4170 3840 4566 3841
rect 4170 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4566 3840
rect 4170 3775 4566 3776
rect 10170 3840 10566 3841
rect 10170 3776 10176 3840
rect 10240 3776 10256 3840
rect 10320 3776 10336 3840
rect 10400 3776 10416 3840
rect 10480 3776 10496 3840
rect 10560 3776 10566 3840
rect 10170 3775 10566 3776
rect 16170 3840 16566 3841
rect 16170 3776 16176 3840
rect 16240 3776 16256 3840
rect 16320 3776 16336 3840
rect 16400 3776 16416 3840
rect 16480 3776 16496 3840
rect 16560 3776 16566 3840
rect 16170 3775 16566 3776
rect 22170 3840 22566 3841
rect 22170 3776 22176 3840
rect 22240 3776 22256 3840
rect 22320 3776 22336 3840
rect 22400 3776 22416 3840
rect 22480 3776 22496 3840
rect 22560 3776 22566 3840
rect 22170 3775 22566 3776
rect 28170 3840 28566 3841
rect 28170 3776 28176 3840
rect 28240 3776 28256 3840
rect 28320 3776 28336 3840
rect 28400 3776 28416 3840
rect 28480 3776 28496 3840
rect 28560 3776 28566 3840
rect 28170 3775 28566 3776
rect 4910 3296 5306 3297
rect 4910 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5306 3296
rect 4910 3231 5306 3232
rect 10910 3296 11306 3297
rect 10910 3232 10916 3296
rect 10980 3232 10996 3296
rect 11060 3232 11076 3296
rect 11140 3232 11156 3296
rect 11220 3232 11236 3296
rect 11300 3232 11306 3296
rect 10910 3231 11306 3232
rect 16910 3296 17306 3297
rect 16910 3232 16916 3296
rect 16980 3232 16996 3296
rect 17060 3232 17076 3296
rect 17140 3232 17156 3296
rect 17220 3232 17236 3296
rect 17300 3232 17306 3296
rect 16910 3231 17306 3232
rect 22910 3296 23306 3297
rect 22910 3232 22916 3296
rect 22980 3232 22996 3296
rect 23060 3232 23076 3296
rect 23140 3232 23156 3296
rect 23220 3232 23236 3296
rect 23300 3232 23306 3296
rect 22910 3231 23306 3232
rect 28910 3296 29306 3297
rect 28910 3232 28916 3296
rect 28980 3232 28996 3296
rect 29060 3232 29076 3296
rect 29140 3232 29156 3296
rect 29220 3232 29236 3296
rect 29300 3232 29306 3296
rect 28910 3231 29306 3232
rect 4170 2752 4566 2753
rect 4170 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4566 2752
rect 4170 2687 4566 2688
rect 10170 2752 10566 2753
rect 10170 2688 10176 2752
rect 10240 2688 10256 2752
rect 10320 2688 10336 2752
rect 10400 2688 10416 2752
rect 10480 2688 10496 2752
rect 10560 2688 10566 2752
rect 10170 2687 10566 2688
rect 16170 2752 16566 2753
rect 16170 2688 16176 2752
rect 16240 2688 16256 2752
rect 16320 2688 16336 2752
rect 16400 2688 16416 2752
rect 16480 2688 16496 2752
rect 16560 2688 16566 2752
rect 16170 2687 16566 2688
rect 22170 2752 22566 2753
rect 22170 2688 22176 2752
rect 22240 2688 22256 2752
rect 22320 2688 22336 2752
rect 22400 2688 22416 2752
rect 22480 2688 22496 2752
rect 22560 2688 22566 2752
rect 22170 2687 22566 2688
rect 28170 2752 28566 2753
rect 28170 2688 28176 2752
rect 28240 2688 28256 2752
rect 28320 2688 28336 2752
rect 28400 2688 28416 2752
rect 28480 2688 28496 2752
rect 28560 2688 28566 2752
rect 28170 2687 28566 2688
rect 4910 2208 5306 2209
rect 4910 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5306 2208
rect 4910 2143 5306 2144
rect 10910 2208 11306 2209
rect 10910 2144 10916 2208
rect 10980 2144 10996 2208
rect 11060 2144 11076 2208
rect 11140 2144 11156 2208
rect 11220 2144 11236 2208
rect 11300 2144 11306 2208
rect 10910 2143 11306 2144
rect 16910 2208 17306 2209
rect 16910 2144 16916 2208
rect 16980 2144 16996 2208
rect 17060 2144 17076 2208
rect 17140 2144 17156 2208
rect 17220 2144 17236 2208
rect 17300 2144 17306 2208
rect 16910 2143 17306 2144
rect 22910 2208 23306 2209
rect 22910 2144 22916 2208
rect 22980 2144 22996 2208
rect 23060 2144 23076 2208
rect 23140 2144 23156 2208
rect 23220 2144 23236 2208
rect 23300 2144 23306 2208
rect 22910 2143 23306 2144
rect 28910 2208 29306 2209
rect 28910 2144 28916 2208
rect 28980 2144 28996 2208
rect 29060 2144 29076 2208
rect 29140 2144 29156 2208
rect 29220 2144 29236 2208
rect 29300 2144 29306 2208
rect 28910 2143 29306 2144
rect 30833 1458 30899 1461
rect 31652 1458 32452 1488
rect 30833 1456 32452 1458
rect 30833 1400 30838 1456
rect 30894 1400 32452 1456
rect 30833 1398 32452 1400
rect 30833 1395 30899 1398
rect 31652 1368 32452 1398
<< via3 >>
rect 4176 32124 4240 32128
rect 4176 32068 4180 32124
rect 4180 32068 4236 32124
rect 4236 32068 4240 32124
rect 4176 32064 4240 32068
rect 4256 32124 4320 32128
rect 4256 32068 4260 32124
rect 4260 32068 4316 32124
rect 4316 32068 4320 32124
rect 4256 32064 4320 32068
rect 4336 32124 4400 32128
rect 4336 32068 4340 32124
rect 4340 32068 4396 32124
rect 4396 32068 4400 32124
rect 4336 32064 4400 32068
rect 4416 32124 4480 32128
rect 4416 32068 4420 32124
rect 4420 32068 4476 32124
rect 4476 32068 4480 32124
rect 4416 32064 4480 32068
rect 4496 32124 4560 32128
rect 4496 32068 4500 32124
rect 4500 32068 4556 32124
rect 4556 32068 4560 32124
rect 4496 32064 4560 32068
rect 10176 32124 10240 32128
rect 10176 32068 10180 32124
rect 10180 32068 10236 32124
rect 10236 32068 10240 32124
rect 10176 32064 10240 32068
rect 10256 32124 10320 32128
rect 10256 32068 10260 32124
rect 10260 32068 10316 32124
rect 10316 32068 10320 32124
rect 10256 32064 10320 32068
rect 10336 32124 10400 32128
rect 10336 32068 10340 32124
rect 10340 32068 10396 32124
rect 10396 32068 10400 32124
rect 10336 32064 10400 32068
rect 10416 32124 10480 32128
rect 10416 32068 10420 32124
rect 10420 32068 10476 32124
rect 10476 32068 10480 32124
rect 10416 32064 10480 32068
rect 10496 32124 10560 32128
rect 10496 32068 10500 32124
rect 10500 32068 10556 32124
rect 10556 32068 10560 32124
rect 10496 32064 10560 32068
rect 16176 32124 16240 32128
rect 16176 32068 16180 32124
rect 16180 32068 16236 32124
rect 16236 32068 16240 32124
rect 16176 32064 16240 32068
rect 16256 32124 16320 32128
rect 16256 32068 16260 32124
rect 16260 32068 16316 32124
rect 16316 32068 16320 32124
rect 16256 32064 16320 32068
rect 16336 32124 16400 32128
rect 16336 32068 16340 32124
rect 16340 32068 16396 32124
rect 16396 32068 16400 32124
rect 16336 32064 16400 32068
rect 16416 32124 16480 32128
rect 16416 32068 16420 32124
rect 16420 32068 16476 32124
rect 16476 32068 16480 32124
rect 16416 32064 16480 32068
rect 16496 32124 16560 32128
rect 16496 32068 16500 32124
rect 16500 32068 16556 32124
rect 16556 32068 16560 32124
rect 16496 32064 16560 32068
rect 22176 32124 22240 32128
rect 22176 32068 22180 32124
rect 22180 32068 22236 32124
rect 22236 32068 22240 32124
rect 22176 32064 22240 32068
rect 22256 32124 22320 32128
rect 22256 32068 22260 32124
rect 22260 32068 22316 32124
rect 22316 32068 22320 32124
rect 22256 32064 22320 32068
rect 22336 32124 22400 32128
rect 22336 32068 22340 32124
rect 22340 32068 22396 32124
rect 22396 32068 22400 32124
rect 22336 32064 22400 32068
rect 22416 32124 22480 32128
rect 22416 32068 22420 32124
rect 22420 32068 22476 32124
rect 22476 32068 22480 32124
rect 22416 32064 22480 32068
rect 22496 32124 22560 32128
rect 22496 32068 22500 32124
rect 22500 32068 22556 32124
rect 22556 32068 22560 32124
rect 22496 32064 22560 32068
rect 28176 32124 28240 32128
rect 28176 32068 28180 32124
rect 28180 32068 28236 32124
rect 28236 32068 28240 32124
rect 28176 32064 28240 32068
rect 28256 32124 28320 32128
rect 28256 32068 28260 32124
rect 28260 32068 28316 32124
rect 28316 32068 28320 32124
rect 28256 32064 28320 32068
rect 28336 32124 28400 32128
rect 28336 32068 28340 32124
rect 28340 32068 28396 32124
rect 28396 32068 28400 32124
rect 28336 32064 28400 32068
rect 28416 32124 28480 32128
rect 28416 32068 28420 32124
rect 28420 32068 28476 32124
rect 28476 32068 28480 32124
rect 28416 32064 28480 32068
rect 28496 32124 28560 32128
rect 28496 32068 28500 32124
rect 28500 32068 28556 32124
rect 28556 32068 28560 32124
rect 28496 32064 28560 32068
rect 24348 31724 24412 31788
rect 4916 31580 4980 31584
rect 4916 31524 4920 31580
rect 4920 31524 4976 31580
rect 4976 31524 4980 31580
rect 4916 31520 4980 31524
rect 4996 31580 5060 31584
rect 4996 31524 5000 31580
rect 5000 31524 5056 31580
rect 5056 31524 5060 31580
rect 4996 31520 5060 31524
rect 5076 31580 5140 31584
rect 5076 31524 5080 31580
rect 5080 31524 5136 31580
rect 5136 31524 5140 31580
rect 5076 31520 5140 31524
rect 5156 31580 5220 31584
rect 5156 31524 5160 31580
rect 5160 31524 5216 31580
rect 5216 31524 5220 31580
rect 5156 31520 5220 31524
rect 5236 31580 5300 31584
rect 5236 31524 5240 31580
rect 5240 31524 5296 31580
rect 5296 31524 5300 31580
rect 5236 31520 5300 31524
rect 10916 31580 10980 31584
rect 10916 31524 10920 31580
rect 10920 31524 10976 31580
rect 10976 31524 10980 31580
rect 10916 31520 10980 31524
rect 10996 31580 11060 31584
rect 10996 31524 11000 31580
rect 11000 31524 11056 31580
rect 11056 31524 11060 31580
rect 10996 31520 11060 31524
rect 11076 31580 11140 31584
rect 11076 31524 11080 31580
rect 11080 31524 11136 31580
rect 11136 31524 11140 31580
rect 11076 31520 11140 31524
rect 11156 31580 11220 31584
rect 11156 31524 11160 31580
rect 11160 31524 11216 31580
rect 11216 31524 11220 31580
rect 11156 31520 11220 31524
rect 11236 31580 11300 31584
rect 11236 31524 11240 31580
rect 11240 31524 11296 31580
rect 11296 31524 11300 31580
rect 11236 31520 11300 31524
rect 16916 31580 16980 31584
rect 16916 31524 16920 31580
rect 16920 31524 16976 31580
rect 16976 31524 16980 31580
rect 16916 31520 16980 31524
rect 16996 31580 17060 31584
rect 16996 31524 17000 31580
rect 17000 31524 17056 31580
rect 17056 31524 17060 31580
rect 16996 31520 17060 31524
rect 17076 31580 17140 31584
rect 17076 31524 17080 31580
rect 17080 31524 17136 31580
rect 17136 31524 17140 31580
rect 17076 31520 17140 31524
rect 17156 31580 17220 31584
rect 17156 31524 17160 31580
rect 17160 31524 17216 31580
rect 17216 31524 17220 31580
rect 17156 31520 17220 31524
rect 17236 31580 17300 31584
rect 17236 31524 17240 31580
rect 17240 31524 17296 31580
rect 17296 31524 17300 31580
rect 17236 31520 17300 31524
rect 22916 31580 22980 31584
rect 22916 31524 22920 31580
rect 22920 31524 22976 31580
rect 22976 31524 22980 31580
rect 22916 31520 22980 31524
rect 22996 31580 23060 31584
rect 22996 31524 23000 31580
rect 23000 31524 23056 31580
rect 23056 31524 23060 31580
rect 22996 31520 23060 31524
rect 23076 31580 23140 31584
rect 23076 31524 23080 31580
rect 23080 31524 23136 31580
rect 23136 31524 23140 31580
rect 23076 31520 23140 31524
rect 23156 31580 23220 31584
rect 23156 31524 23160 31580
rect 23160 31524 23216 31580
rect 23216 31524 23220 31580
rect 23156 31520 23220 31524
rect 23236 31580 23300 31584
rect 23236 31524 23240 31580
rect 23240 31524 23296 31580
rect 23296 31524 23300 31580
rect 23236 31520 23300 31524
rect 28916 31580 28980 31584
rect 28916 31524 28920 31580
rect 28920 31524 28976 31580
rect 28976 31524 28980 31580
rect 28916 31520 28980 31524
rect 28996 31580 29060 31584
rect 28996 31524 29000 31580
rect 29000 31524 29056 31580
rect 29056 31524 29060 31580
rect 28996 31520 29060 31524
rect 29076 31580 29140 31584
rect 29076 31524 29080 31580
rect 29080 31524 29136 31580
rect 29136 31524 29140 31580
rect 29076 31520 29140 31524
rect 29156 31580 29220 31584
rect 29156 31524 29160 31580
rect 29160 31524 29216 31580
rect 29216 31524 29220 31580
rect 29156 31520 29220 31524
rect 29236 31580 29300 31584
rect 29236 31524 29240 31580
rect 29240 31524 29296 31580
rect 29296 31524 29300 31580
rect 29236 31520 29300 31524
rect 27844 31316 27908 31380
rect 4176 31036 4240 31040
rect 4176 30980 4180 31036
rect 4180 30980 4236 31036
rect 4236 30980 4240 31036
rect 4176 30976 4240 30980
rect 4256 31036 4320 31040
rect 4256 30980 4260 31036
rect 4260 30980 4316 31036
rect 4316 30980 4320 31036
rect 4256 30976 4320 30980
rect 4336 31036 4400 31040
rect 4336 30980 4340 31036
rect 4340 30980 4396 31036
rect 4396 30980 4400 31036
rect 4336 30976 4400 30980
rect 4416 31036 4480 31040
rect 4416 30980 4420 31036
rect 4420 30980 4476 31036
rect 4476 30980 4480 31036
rect 4416 30976 4480 30980
rect 4496 31036 4560 31040
rect 4496 30980 4500 31036
rect 4500 30980 4556 31036
rect 4556 30980 4560 31036
rect 4496 30976 4560 30980
rect 10176 31036 10240 31040
rect 10176 30980 10180 31036
rect 10180 30980 10236 31036
rect 10236 30980 10240 31036
rect 10176 30976 10240 30980
rect 10256 31036 10320 31040
rect 10256 30980 10260 31036
rect 10260 30980 10316 31036
rect 10316 30980 10320 31036
rect 10256 30976 10320 30980
rect 10336 31036 10400 31040
rect 10336 30980 10340 31036
rect 10340 30980 10396 31036
rect 10396 30980 10400 31036
rect 10336 30976 10400 30980
rect 10416 31036 10480 31040
rect 10416 30980 10420 31036
rect 10420 30980 10476 31036
rect 10476 30980 10480 31036
rect 10416 30976 10480 30980
rect 10496 31036 10560 31040
rect 10496 30980 10500 31036
rect 10500 30980 10556 31036
rect 10556 30980 10560 31036
rect 10496 30976 10560 30980
rect 16176 31036 16240 31040
rect 16176 30980 16180 31036
rect 16180 30980 16236 31036
rect 16236 30980 16240 31036
rect 16176 30976 16240 30980
rect 16256 31036 16320 31040
rect 16256 30980 16260 31036
rect 16260 30980 16316 31036
rect 16316 30980 16320 31036
rect 16256 30976 16320 30980
rect 16336 31036 16400 31040
rect 16336 30980 16340 31036
rect 16340 30980 16396 31036
rect 16396 30980 16400 31036
rect 16336 30976 16400 30980
rect 16416 31036 16480 31040
rect 16416 30980 16420 31036
rect 16420 30980 16476 31036
rect 16476 30980 16480 31036
rect 16416 30976 16480 30980
rect 16496 31036 16560 31040
rect 16496 30980 16500 31036
rect 16500 30980 16556 31036
rect 16556 30980 16560 31036
rect 16496 30976 16560 30980
rect 22176 31036 22240 31040
rect 22176 30980 22180 31036
rect 22180 30980 22236 31036
rect 22236 30980 22240 31036
rect 22176 30976 22240 30980
rect 22256 31036 22320 31040
rect 22256 30980 22260 31036
rect 22260 30980 22316 31036
rect 22316 30980 22320 31036
rect 22256 30976 22320 30980
rect 22336 31036 22400 31040
rect 22336 30980 22340 31036
rect 22340 30980 22396 31036
rect 22396 30980 22400 31036
rect 22336 30976 22400 30980
rect 22416 31036 22480 31040
rect 22416 30980 22420 31036
rect 22420 30980 22476 31036
rect 22476 30980 22480 31036
rect 22416 30976 22480 30980
rect 22496 31036 22560 31040
rect 22496 30980 22500 31036
rect 22500 30980 22556 31036
rect 22556 30980 22560 31036
rect 22496 30976 22560 30980
rect 28176 31036 28240 31040
rect 28176 30980 28180 31036
rect 28180 30980 28236 31036
rect 28236 30980 28240 31036
rect 28176 30976 28240 30980
rect 28256 31036 28320 31040
rect 28256 30980 28260 31036
rect 28260 30980 28316 31036
rect 28316 30980 28320 31036
rect 28256 30976 28320 30980
rect 28336 31036 28400 31040
rect 28336 30980 28340 31036
rect 28340 30980 28396 31036
rect 28396 30980 28400 31036
rect 28336 30976 28400 30980
rect 28416 31036 28480 31040
rect 28416 30980 28420 31036
rect 28420 30980 28476 31036
rect 28476 30980 28480 31036
rect 28416 30976 28480 30980
rect 28496 31036 28560 31040
rect 28496 30980 28500 31036
rect 28500 30980 28556 31036
rect 28556 30980 28560 31036
rect 28496 30976 28560 30980
rect 4916 30492 4980 30496
rect 4916 30436 4920 30492
rect 4920 30436 4976 30492
rect 4976 30436 4980 30492
rect 4916 30432 4980 30436
rect 4996 30492 5060 30496
rect 4996 30436 5000 30492
rect 5000 30436 5056 30492
rect 5056 30436 5060 30492
rect 4996 30432 5060 30436
rect 5076 30492 5140 30496
rect 5076 30436 5080 30492
rect 5080 30436 5136 30492
rect 5136 30436 5140 30492
rect 5076 30432 5140 30436
rect 5156 30492 5220 30496
rect 5156 30436 5160 30492
rect 5160 30436 5216 30492
rect 5216 30436 5220 30492
rect 5156 30432 5220 30436
rect 5236 30492 5300 30496
rect 5236 30436 5240 30492
rect 5240 30436 5296 30492
rect 5296 30436 5300 30492
rect 5236 30432 5300 30436
rect 10916 30492 10980 30496
rect 10916 30436 10920 30492
rect 10920 30436 10976 30492
rect 10976 30436 10980 30492
rect 10916 30432 10980 30436
rect 10996 30492 11060 30496
rect 10996 30436 11000 30492
rect 11000 30436 11056 30492
rect 11056 30436 11060 30492
rect 10996 30432 11060 30436
rect 11076 30492 11140 30496
rect 11076 30436 11080 30492
rect 11080 30436 11136 30492
rect 11136 30436 11140 30492
rect 11076 30432 11140 30436
rect 11156 30492 11220 30496
rect 11156 30436 11160 30492
rect 11160 30436 11216 30492
rect 11216 30436 11220 30492
rect 11156 30432 11220 30436
rect 11236 30492 11300 30496
rect 11236 30436 11240 30492
rect 11240 30436 11296 30492
rect 11296 30436 11300 30492
rect 11236 30432 11300 30436
rect 16916 30492 16980 30496
rect 16916 30436 16920 30492
rect 16920 30436 16976 30492
rect 16976 30436 16980 30492
rect 16916 30432 16980 30436
rect 16996 30492 17060 30496
rect 16996 30436 17000 30492
rect 17000 30436 17056 30492
rect 17056 30436 17060 30492
rect 16996 30432 17060 30436
rect 17076 30492 17140 30496
rect 17076 30436 17080 30492
rect 17080 30436 17136 30492
rect 17136 30436 17140 30492
rect 17076 30432 17140 30436
rect 17156 30492 17220 30496
rect 17156 30436 17160 30492
rect 17160 30436 17216 30492
rect 17216 30436 17220 30492
rect 17156 30432 17220 30436
rect 17236 30492 17300 30496
rect 17236 30436 17240 30492
rect 17240 30436 17296 30492
rect 17296 30436 17300 30492
rect 17236 30432 17300 30436
rect 22916 30492 22980 30496
rect 22916 30436 22920 30492
rect 22920 30436 22976 30492
rect 22976 30436 22980 30492
rect 22916 30432 22980 30436
rect 22996 30492 23060 30496
rect 22996 30436 23000 30492
rect 23000 30436 23056 30492
rect 23056 30436 23060 30492
rect 22996 30432 23060 30436
rect 23076 30492 23140 30496
rect 23076 30436 23080 30492
rect 23080 30436 23136 30492
rect 23136 30436 23140 30492
rect 23076 30432 23140 30436
rect 23156 30492 23220 30496
rect 23156 30436 23160 30492
rect 23160 30436 23216 30492
rect 23216 30436 23220 30492
rect 23156 30432 23220 30436
rect 23236 30492 23300 30496
rect 23236 30436 23240 30492
rect 23240 30436 23296 30492
rect 23296 30436 23300 30492
rect 23236 30432 23300 30436
rect 28916 30492 28980 30496
rect 28916 30436 28920 30492
rect 28920 30436 28976 30492
rect 28976 30436 28980 30492
rect 28916 30432 28980 30436
rect 28996 30492 29060 30496
rect 28996 30436 29000 30492
rect 29000 30436 29056 30492
rect 29056 30436 29060 30492
rect 28996 30432 29060 30436
rect 29076 30492 29140 30496
rect 29076 30436 29080 30492
rect 29080 30436 29136 30492
rect 29136 30436 29140 30492
rect 29076 30432 29140 30436
rect 29156 30492 29220 30496
rect 29156 30436 29160 30492
rect 29160 30436 29216 30492
rect 29216 30436 29220 30492
rect 29156 30432 29220 30436
rect 29236 30492 29300 30496
rect 29236 30436 29240 30492
rect 29240 30436 29296 30492
rect 29296 30436 29300 30492
rect 29236 30432 29300 30436
rect 4176 29948 4240 29952
rect 4176 29892 4180 29948
rect 4180 29892 4236 29948
rect 4236 29892 4240 29948
rect 4176 29888 4240 29892
rect 4256 29948 4320 29952
rect 4256 29892 4260 29948
rect 4260 29892 4316 29948
rect 4316 29892 4320 29948
rect 4256 29888 4320 29892
rect 4336 29948 4400 29952
rect 4336 29892 4340 29948
rect 4340 29892 4396 29948
rect 4396 29892 4400 29948
rect 4336 29888 4400 29892
rect 4416 29948 4480 29952
rect 4416 29892 4420 29948
rect 4420 29892 4476 29948
rect 4476 29892 4480 29948
rect 4416 29888 4480 29892
rect 4496 29948 4560 29952
rect 4496 29892 4500 29948
rect 4500 29892 4556 29948
rect 4556 29892 4560 29948
rect 4496 29888 4560 29892
rect 10176 29948 10240 29952
rect 10176 29892 10180 29948
rect 10180 29892 10236 29948
rect 10236 29892 10240 29948
rect 10176 29888 10240 29892
rect 10256 29948 10320 29952
rect 10256 29892 10260 29948
rect 10260 29892 10316 29948
rect 10316 29892 10320 29948
rect 10256 29888 10320 29892
rect 10336 29948 10400 29952
rect 10336 29892 10340 29948
rect 10340 29892 10396 29948
rect 10396 29892 10400 29948
rect 10336 29888 10400 29892
rect 10416 29948 10480 29952
rect 10416 29892 10420 29948
rect 10420 29892 10476 29948
rect 10476 29892 10480 29948
rect 10416 29888 10480 29892
rect 10496 29948 10560 29952
rect 10496 29892 10500 29948
rect 10500 29892 10556 29948
rect 10556 29892 10560 29948
rect 10496 29888 10560 29892
rect 16176 29948 16240 29952
rect 16176 29892 16180 29948
rect 16180 29892 16236 29948
rect 16236 29892 16240 29948
rect 16176 29888 16240 29892
rect 16256 29948 16320 29952
rect 16256 29892 16260 29948
rect 16260 29892 16316 29948
rect 16316 29892 16320 29948
rect 16256 29888 16320 29892
rect 16336 29948 16400 29952
rect 16336 29892 16340 29948
rect 16340 29892 16396 29948
rect 16396 29892 16400 29948
rect 16336 29888 16400 29892
rect 16416 29948 16480 29952
rect 16416 29892 16420 29948
rect 16420 29892 16476 29948
rect 16476 29892 16480 29948
rect 16416 29888 16480 29892
rect 16496 29948 16560 29952
rect 16496 29892 16500 29948
rect 16500 29892 16556 29948
rect 16556 29892 16560 29948
rect 16496 29888 16560 29892
rect 22176 29948 22240 29952
rect 22176 29892 22180 29948
rect 22180 29892 22236 29948
rect 22236 29892 22240 29948
rect 22176 29888 22240 29892
rect 22256 29948 22320 29952
rect 22256 29892 22260 29948
rect 22260 29892 22316 29948
rect 22316 29892 22320 29948
rect 22256 29888 22320 29892
rect 22336 29948 22400 29952
rect 22336 29892 22340 29948
rect 22340 29892 22396 29948
rect 22396 29892 22400 29948
rect 22336 29888 22400 29892
rect 22416 29948 22480 29952
rect 22416 29892 22420 29948
rect 22420 29892 22476 29948
rect 22476 29892 22480 29948
rect 22416 29888 22480 29892
rect 22496 29948 22560 29952
rect 22496 29892 22500 29948
rect 22500 29892 22556 29948
rect 22556 29892 22560 29948
rect 22496 29888 22560 29892
rect 28176 29948 28240 29952
rect 28176 29892 28180 29948
rect 28180 29892 28236 29948
rect 28236 29892 28240 29948
rect 28176 29888 28240 29892
rect 28256 29948 28320 29952
rect 28256 29892 28260 29948
rect 28260 29892 28316 29948
rect 28316 29892 28320 29948
rect 28256 29888 28320 29892
rect 28336 29948 28400 29952
rect 28336 29892 28340 29948
rect 28340 29892 28396 29948
rect 28396 29892 28400 29948
rect 28336 29888 28400 29892
rect 28416 29948 28480 29952
rect 28416 29892 28420 29948
rect 28420 29892 28476 29948
rect 28476 29892 28480 29948
rect 28416 29888 28480 29892
rect 28496 29948 28560 29952
rect 28496 29892 28500 29948
rect 28500 29892 28556 29948
rect 28556 29892 28560 29948
rect 28496 29888 28560 29892
rect 4916 29404 4980 29408
rect 4916 29348 4920 29404
rect 4920 29348 4976 29404
rect 4976 29348 4980 29404
rect 4916 29344 4980 29348
rect 4996 29404 5060 29408
rect 4996 29348 5000 29404
rect 5000 29348 5056 29404
rect 5056 29348 5060 29404
rect 4996 29344 5060 29348
rect 5076 29404 5140 29408
rect 5076 29348 5080 29404
rect 5080 29348 5136 29404
rect 5136 29348 5140 29404
rect 5076 29344 5140 29348
rect 5156 29404 5220 29408
rect 5156 29348 5160 29404
rect 5160 29348 5216 29404
rect 5216 29348 5220 29404
rect 5156 29344 5220 29348
rect 5236 29404 5300 29408
rect 5236 29348 5240 29404
rect 5240 29348 5296 29404
rect 5296 29348 5300 29404
rect 5236 29344 5300 29348
rect 10916 29404 10980 29408
rect 10916 29348 10920 29404
rect 10920 29348 10976 29404
rect 10976 29348 10980 29404
rect 10916 29344 10980 29348
rect 10996 29404 11060 29408
rect 10996 29348 11000 29404
rect 11000 29348 11056 29404
rect 11056 29348 11060 29404
rect 10996 29344 11060 29348
rect 11076 29404 11140 29408
rect 11076 29348 11080 29404
rect 11080 29348 11136 29404
rect 11136 29348 11140 29404
rect 11076 29344 11140 29348
rect 11156 29404 11220 29408
rect 11156 29348 11160 29404
rect 11160 29348 11216 29404
rect 11216 29348 11220 29404
rect 11156 29344 11220 29348
rect 11236 29404 11300 29408
rect 11236 29348 11240 29404
rect 11240 29348 11296 29404
rect 11296 29348 11300 29404
rect 11236 29344 11300 29348
rect 16916 29404 16980 29408
rect 16916 29348 16920 29404
rect 16920 29348 16976 29404
rect 16976 29348 16980 29404
rect 16916 29344 16980 29348
rect 16996 29404 17060 29408
rect 16996 29348 17000 29404
rect 17000 29348 17056 29404
rect 17056 29348 17060 29404
rect 16996 29344 17060 29348
rect 17076 29404 17140 29408
rect 17076 29348 17080 29404
rect 17080 29348 17136 29404
rect 17136 29348 17140 29404
rect 17076 29344 17140 29348
rect 17156 29404 17220 29408
rect 17156 29348 17160 29404
rect 17160 29348 17216 29404
rect 17216 29348 17220 29404
rect 17156 29344 17220 29348
rect 17236 29404 17300 29408
rect 17236 29348 17240 29404
rect 17240 29348 17296 29404
rect 17296 29348 17300 29404
rect 17236 29344 17300 29348
rect 22916 29404 22980 29408
rect 22916 29348 22920 29404
rect 22920 29348 22976 29404
rect 22976 29348 22980 29404
rect 22916 29344 22980 29348
rect 22996 29404 23060 29408
rect 22996 29348 23000 29404
rect 23000 29348 23056 29404
rect 23056 29348 23060 29404
rect 22996 29344 23060 29348
rect 23076 29404 23140 29408
rect 23076 29348 23080 29404
rect 23080 29348 23136 29404
rect 23136 29348 23140 29404
rect 23076 29344 23140 29348
rect 23156 29404 23220 29408
rect 23156 29348 23160 29404
rect 23160 29348 23216 29404
rect 23216 29348 23220 29404
rect 23156 29344 23220 29348
rect 23236 29404 23300 29408
rect 23236 29348 23240 29404
rect 23240 29348 23296 29404
rect 23296 29348 23300 29404
rect 23236 29344 23300 29348
rect 28916 29404 28980 29408
rect 28916 29348 28920 29404
rect 28920 29348 28976 29404
rect 28976 29348 28980 29404
rect 28916 29344 28980 29348
rect 28996 29404 29060 29408
rect 28996 29348 29000 29404
rect 29000 29348 29056 29404
rect 29056 29348 29060 29404
rect 28996 29344 29060 29348
rect 29076 29404 29140 29408
rect 29076 29348 29080 29404
rect 29080 29348 29136 29404
rect 29136 29348 29140 29404
rect 29076 29344 29140 29348
rect 29156 29404 29220 29408
rect 29156 29348 29160 29404
rect 29160 29348 29216 29404
rect 29216 29348 29220 29404
rect 29156 29344 29220 29348
rect 29236 29404 29300 29408
rect 29236 29348 29240 29404
rect 29240 29348 29296 29404
rect 29296 29348 29300 29404
rect 29236 29344 29300 29348
rect 4176 28860 4240 28864
rect 4176 28804 4180 28860
rect 4180 28804 4236 28860
rect 4236 28804 4240 28860
rect 4176 28800 4240 28804
rect 4256 28860 4320 28864
rect 4256 28804 4260 28860
rect 4260 28804 4316 28860
rect 4316 28804 4320 28860
rect 4256 28800 4320 28804
rect 4336 28860 4400 28864
rect 4336 28804 4340 28860
rect 4340 28804 4396 28860
rect 4396 28804 4400 28860
rect 4336 28800 4400 28804
rect 4416 28860 4480 28864
rect 4416 28804 4420 28860
rect 4420 28804 4476 28860
rect 4476 28804 4480 28860
rect 4416 28800 4480 28804
rect 4496 28860 4560 28864
rect 4496 28804 4500 28860
rect 4500 28804 4556 28860
rect 4556 28804 4560 28860
rect 4496 28800 4560 28804
rect 10176 28860 10240 28864
rect 10176 28804 10180 28860
rect 10180 28804 10236 28860
rect 10236 28804 10240 28860
rect 10176 28800 10240 28804
rect 10256 28860 10320 28864
rect 10256 28804 10260 28860
rect 10260 28804 10316 28860
rect 10316 28804 10320 28860
rect 10256 28800 10320 28804
rect 10336 28860 10400 28864
rect 10336 28804 10340 28860
rect 10340 28804 10396 28860
rect 10396 28804 10400 28860
rect 10336 28800 10400 28804
rect 10416 28860 10480 28864
rect 10416 28804 10420 28860
rect 10420 28804 10476 28860
rect 10476 28804 10480 28860
rect 10416 28800 10480 28804
rect 10496 28860 10560 28864
rect 10496 28804 10500 28860
rect 10500 28804 10556 28860
rect 10556 28804 10560 28860
rect 10496 28800 10560 28804
rect 16176 28860 16240 28864
rect 16176 28804 16180 28860
rect 16180 28804 16236 28860
rect 16236 28804 16240 28860
rect 16176 28800 16240 28804
rect 16256 28860 16320 28864
rect 16256 28804 16260 28860
rect 16260 28804 16316 28860
rect 16316 28804 16320 28860
rect 16256 28800 16320 28804
rect 16336 28860 16400 28864
rect 16336 28804 16340 28860
rect 16340 28804 16396 28860
rect 16396 28804 16400 28860
rect 16336 28800 16400 28804
rect 16416 28860 16480 28864
rect 16416 28804 16420 28860
rect 16420 28804 16476 28860
rect 16476 28804 16480 28860
rect 16416 28800 16480 28804
rect 16496 28860 16560 28864
rect 16496 28804 16500 28860
rect 16500 28804 16556 28860
rect 16556 28804 16560 28860
rect 16496 28800 16560 28804
rect 22176 28860 22240 28864
rect 22176 28804 22180 28860
rect 22180 28804 22236 28860
rect 22236 28804 22240 28860
rect 22176 28800 22240 28804
rect 22256 28860 22320 28864
rect 22256 28804 22260 28860
rect 22260 28804 22316 28860
rect 22316 28804 22320 28860
rect 22256 28800 22320 28804
rect 22336 28860 22400 28864
rect 22336 28804 22340 28860
rect 22340 28804 22396 28860
rect 22396 28804 22400 28860
rect 22336 28800 22400 28804
rect 22416 28860 22480 28864
rect 22416 28804 22420 28860
rect 22420 28804 22476 28860
rect 22476 28804 22480 28860
rect 22416 28800 22480 28804
rect 22496 28860 22560 28864
rect 22496 28804 22500 28860
rect 22500 28804 22556 28860
rect 22556 28804 22560 28860
rect 22496 28800 22560 28804
rect 28176 28860 28240 28864
rect 28176 28804 28180 28860
rect 28180 28804 28236 28860
rect 28236 28804 28240 28860
rect 28176 28800 28240 28804
rect 28256 28860 28320 28864
rect 28256 28804 28260 28860
rect 28260 28804 28316 28860
rect 28316 28804 28320 28860
rect 28256 28800 28320 28804
rect 28336 28860 28400 28864
rect 28336 28804 28340 28860
rect 28340 28804 28396 28860
rect 28396 28804 28400 28860
rect 28336 28800 28400 28804
rect 28416 28860 28480 28864
rect 28416 28804 28420 28860
rect 28420 28804 28476 28860
rect 28476 28804 28480 28860
rect 28416 28800 28480 28804
rect 28496 28860 28560 28864
rect 28496 28804 28500 28860
rect 28500 28804 28556 28860
rect 28556 28804 28560 28860
rect 28496 28800 28560 28804
rect 4916 28316 4980 28320
rect 4916 28260 4920 28316
rect 4920 28260 4976 28316
rect 4976 28260 4980 28316
rect 4916 28256 4980 28260
rect 4996 28316 5060 28320
rect 4996 28260 5000 28316
rect 5000 28260 5056 28316
rect 5056 28260 5060 28316
rect 4996 28256 5060 28260
rect 5076 28316 5140 28320
rect 5076 28260 5080 28316
rect 5080 28260 5136 28316
rect 5136 28260 5140 28316
rect 5076 28256 5140 28260
rect 5156 28316 5220 28320
rect 5156 28260 5160 28316
rect 5160 28260 5216 28316
rect 5216 28260 5220 28316
rect 5156 28256 5220 28260
rect 5236 28316 5300 28320
rect 5236 28260 5240 28316
rect 5240 28260 5296 28316
rect 5296 28260 5300 28316
rect 5236 28256 5300 28260
rect 10916 28316 10980 28320
rect 10916 28260 10920 28316
rect 10920 28260 10976 28316
rect 10976 28260 10980 28316
rect 10916 28256 10980 28260
rect 10996 28316 11060 28320
rect 10996 28260 11000 28316
rect 11000 28260 11056 28316
rect 11056 28260 11060 28316
rect 10996 28256 11060 28260
rect 11076 28316 11140 28320
rect 11076 28260 11080 28316
rect 11080 28260 11136 28316
rect 11136 28260 11140 28316
rect 11076 28256 11140 28260
rect 11156 28316 11220 28320
rect 11156 28260 11160 28316
rect 11160 28260 11216 28316
rect 11216 28260 11220 28316
rect 11156 28256 11220 28260
rect 11236 28316 11300 28320
rect 11236 28260 11240 28316
rect 11240 28260 11296 28316
rect 11296 28260 11300 28316
rect 11236 28256 11300 28260
rect 16916 28316 16980 28320
rect 16916 28260 16920 28316
rect 16920 28260 16976 28316
rect 16976 28260 16980 28316
rect 16916 28256 16980 28260
rect 16996 28316 17060 28320
rect 16996 28260 17000 28316
rect 17000 28260 17056 28316
rect 17056 28260 17060 28316
rect 16996 28256 17060 28260
rect 17076 28316 17140 28320
rect 17076 28260 17080 28316
rect 17080 28260 17136 28316
rect 17136 28260 17140 28316
rect 17076 28256 17140 28260
rect 17156 28316 17220 28320
rect 17156 28260 17160 28316
rect 17160 28260 17216 28316
rect 17216 28260 17220 28316
rect 17156 28256 17220 28260
rect 17236 28316 17300 28320
rect 17236 28260 17240 28316
rect 17240 28260 17296 28316
rect 17296 28260 17300 28316
rect 17236 28256 17300 28260
rect 22916 28316 22980 28320
rect 22916 28260 22920 28316
rect 22920 28260 22976 28316
rect 22976 28260 22980 28316
rect 22916 28256 22980 28260
rect 22996 28316 23060 28320
rect 22996 28260 23000 28316
rect 23000 28260 23056 28316
rect 23056 28260 23060 28316
rect 22996 28256 23060 28260
rect 23076 28316 23140 28320
rect 23076 28260 23080 28316
rect 23080 28260 23136 28316
rect 23136 28260 23140 28316
rect 23076 28256 23140 28260
rect 23156 28316 23220 28320
rect 23156 28260 23160 28316
rect 23160 28260 23216 28316
rect 23216 28260 23220 28316
rect 23156 28256 23220 28260
rect 23236 28316 23300 28320
rect 23236 28260 23240 28316
rect 23240 28260 23296 28316
rect 23296 28260 23300 28316
rect 23236 28256 23300 28260
rect 28916 28316 28980 28320
rect 28916 28260 28920 28316
rect 28920 28260 28976 28316
rect 28976 28260 28980 28316
rect 28916 28256 28980 28260
rect 28996 28316 29060 28320
rect 28996 28260 29000 28316
rect 29000 28260 29056 28316
rect 29056 28260 29060 28316
rect 28996 28256 29060 28260
rect 29076 28316 29140 28320
rect 29076 28260 29080 28316
rect 29080 28260 29136 28316
rect 29136 28260 29140 28316
rect 29076 28256 29140 28260
rect 29156 28316 29220 28320
rect 29156 28260 29160 28316
rect 29160 28260 29216 28316
rect 29216 28260 29220 28316
rect 29156 28256 29220 28260
rect 29236 28316 29300 28320
rect 29236 28260 29240 28316
rect 29240 28260 29296 28316
rect 29296 28260 29300 28316
rect 29236 28256 29300 28260
rect 4176 27772 4240 27776
rect 4176 27716 4180 27772
rect 4180 27716 4236 27772
rect 4236 27716 4240 27772
rect 4176 27712 4240 27716
rect 4256 27772 4320 27776
rect 4256 27716 4260 27772
rect 4260 27716 4316 27772
rect 4316 27716 4320 27772
rect 4256 27712 4320 27716
rect 4336 27772 4400 27776
rect 4336 27716 4340 27772
rect 4340 27716 4396 27772
rect 4396 27716 4400 27772
rect 4336 27712 4400 27716
rect 4416 27772 4480 27776
rect 4416 27716 4420 27772
rect 4420 27716 4476 27772
rect 4476 27716 4480 27772
rect 4416 27712 4480 27716
rect 4496 27772 4560 27776
rect 4496 27716 4500 27772
rect 4500 27716 4556 27772
rect 4556 27716 4560 27772
rect 4496 27712 4560 27716
rect 10176 27772 10240 27776
rect 10176 27716 10180 27772
rect 10180 27716 10236 27772
rect 10236 27716 10240 27772
rect 10176 27712 10240 27716
rect 10256 27772 10320 27776
rect 10256 27716 10260 27772
rect 10260 27716 10316 27772
rect 10316 27716 10320 27772
rect 10256 27712 10320 27716
rect 10336 27772 10400 27776
rect 10336 27716 10340 27772
rect 10340 27716 10396 27772
rect 10396 27716 10400 27772
rect 10336 27712 10400 27716
rect 10416 27772 10480 27776
rect 10416 27716 10420 27772
rect 10420 27716 10476 27772
rect 10476 27716 10480 27772
rect 10416 27712 10480 27716
rect 10496 27772 10560 27776
rect 10496 27716 10500 27772
rect 10500 27716 10556 27772
rect 10556 27716 10560 27772
rect 10496 27712 10560 27716
rect 16176 27772 16240 27776
rect 16176 27716 16180 27772
rect 16180 27716 16236 27772
rect 16236 27716 16240 27772
rect 16176 27712 16240 27716
rect 16256 27772 16320 27776
rect 16256 27716 16260 27772
rect 16260 27716 16316 27772
rect 16316 27716 16320 27772
rect 16256 27712 16320 27716
rect 16336 27772 16400 27776
rect 16336 27716 16340 27772
rect 16340 27716 16396 27772
rect 16396 27716 16400 27772
rect 16336 27712 16400 27716
rect 16416 27772 16480 27776
rect 16416 27716 16420 27772
rect 16420 27716 16476 27772
rect 16476 27716 16480 27772
rect 16416 27712 16480 27716
rect 16496 27772 16560 27776
rect 16496 27716 16500 27772
rect 16500 27716 16556 27772
rect 16556 27716 16560 27772
rect 16496 27712 16560 27716
rect 22176 27772 22240 27776
rect 22176 27716 22180 27772
rect 22180 27716 22236 27772
rect 22236 27716 22240 27772
rect 22176 27712 22240 27716
rect 22256 27772 22320 27776
rect 22256 27716 22260 27772
rect 22260 27716 22316 27772
rect 22316 27716 22320 27772
rect 22256 27712 22320 27716
rect 22336 27772 22400 27776
rect 22336 27716 22340 27772
rect 22340 27716 22396 27772
rect 22396 27716 22400 27772
rect 22336 27712 22400 27716
rect 22416 27772 22480 27776
rect 22416 27716 22420 27772
rect 22420 27716 22476 27772
rect 22476 27716 22480 27772
rect 22416 27712 22480 27716
rect 22496 27772 22560 27776
rect 22496 27716 22500 27772
rect 22500 27716 22556 27772
rect 22556 27716 22560 27772
rect 22496 27712 22560 27716
rect 28176 27772 28240 27776
rect 28176 27716 28180 27772
rect 28180 27716 28236 27772
rect 28236 27716 28240 27772
rect 28176 27712 28240 27716
rect 28256 27772 28320 27776
rect 28256 27716 28260 27772
rect 28260 27716 28316 27772
rect 28316 27716 28320 27772
rect 28256 27712 28320 27716
rect 28336 27772 28400 27776
rect 28336 27716 28340 27772
rect 28340 27716 28396 27772
rect 28396 27716 28400 27772
rect 28336 27712 28400 27716
rect 28416 27772 28480 27776
rect 28416 27716 28420 27772
rect 28420 27716 28476 27772
rect 28476 27716 28480 27772
rect 28416 27712 28480 27716
rect 28496 27772 28560 27776
rect 28496 27716 28500 27772
rect 28500 27716 28556 27772
rect 28556 27716 28560 27772
rect 28496 27712 28560 27716
rect 24532 27644 24596 27708
rect 4916 27228 4980 27232
rect 4916 27172 4920 27228
rect 4920 27172 4976 27228
rect 4976 27172 4980 27228
rect 4916 27168 4980 27172
rect 4996 27228 5060 27232
rect 4996 27172 5000 27228
rect 5000 27172 5056 27228
rect 5056 27172 5060 27228
rect 4996 27168 5060 27172
rect 5076 27228 5140 27232
rect 5076 27172 5080 27228
rect 5080 27172 5136 27228
rect 5136 27172 5140 27228
rect 5076 27168 5140 27172
rect 5156 27228 5220 27232
rect 5156 27172 5160 27228
rect 5160 27172 5216 27228
rect 5216 27172 5220 27228
rect 5156 27168 5220 27172
rect 5236 27228 5300 27232
rect 5236 27172 5240 27228
rect 5240 27172 5296 27228
rect 5296 27172 5300 27228
rect 5236 27168 5300 27172
rect 10916 27228 10980 27232
rect 10916 27172 10920 27228
rect 10920 27172 10976 27228
rect 10976 27172 10980 27228
rect 10916 27168 10980 27172
rect 10996 27228 11060 27232
rect 10996 27172 11000 27228
rect 11000 27172 11056 27228
rect 11056 27172 11060 27228
rect 10996 27168 11060 27172
rect 11076 27228 11140 27232
rect 11076 27172 11080 27228
rect 11080 27172 11136 27228
rect 11136 27172 11140 27228
rect 11076 27168 11140 27172
rect 11156 27228 11220 27232
rect 11156 27172 11160 27228
rect 11160 27172 11216 27228
rect 11216 27172 11220 27228
rect 11156 27168 11220 27172
rect 11236 27228 11300 27232
rect 11236 27172 11240 27228
rect 11240 27172 11296 27228
rect 11296 27172 11300 27228
rect 11236 27168 11300 27172
rect 16916 27228 16980 27232
rect 16916 27172 16920 27228
rect 16920 27172 16976 27228
rect 16976 27172 16980 27228
rect 16916 27168 16980 27172
rect 16996 27228 17060 27232
rect 16996 27172 17000 27228
rect 17000 27172 17056 27228
rect 17056 27172 17060 27228
rect 16996 27168 17060 27172
rect 17076 27228 17140 27232
rect 17076 27172 17080 27228
rect 17080 27172 17136 27228
rect 17136 27172 17140 27228
rect 17076 27168 17140 27172
rect 17156 27228 17220 27232
rect 17156 27172 17160 27228
rect 17160 27172 17216 27228
rect 17216 27172 17220 27228
rect 17156 27168 17220 27172
rect 17236 27228 17300 27232
rect 17236 27172 17240 27228
rect 17240 27172 17296 27228
rect 17296 27172 17300 27228
rect 17236 27168 17300 27172
rect 22916 27228 22980 27232
rect 22916 27172 22920 27228
rect 22920 27172 22976 27228
rect 22976 27172 22980 27228
rect 22916 27168 22980 27172
rect 22996 27228 23060 27232
rect 22996 27172 23000 27228
rect 23000 27172 23056 27228
rect 23056 27172 23060 27228
rect 22996 27168 23060 27172
rect 23076 27228 23140 27232
rect 23076 27172 23080 27228
rect 23080 27172 23136 27228
rect 23136 27172 23140 27228
rect 23076 27168 23140 27172
rect 23156 27228 23220 27232
rect 23156 27172 23160 27228
rect 23160 27172 23216 27228
rect 23216 27172 23220 27228
rect 23156 27168 23220 27172
rect 23236 27228 23300 27232
rect 23236 27172 23240 27228
rect 23240 27172 23296 27228
rect 23296 27172 23300 27228
rect 23236 27168 23300 27172
rect 28916 27228 28980 27232
rect 28916 27172 28920 27228
rect 28920 27172 28976 27228
rect 28976 27172 28980 27228
rect 28916 27168 28980 27172
rect 28996 27228 29060 27232
rect 28996 27172 29000 27228
rect 29000 27172 29056 27228
rect 29056 27172 29060 27228
rect 28996 27168 29060 27172
rect 29076 27228 29140 27232
rect 29076 27172 29080 27228
rect 29080 27172 29136 27228
rect 29136 27172 29140 27228
rect 29076 27168 29140 27172
rect 29156 27228 29220 27232
rect 29156 27172 29160 27228
rect 29160 27172 29216 27228
rect 29216 27172 29220 27228
rect 29156 27168 29220 27172
rect 29236 27228 29300 27232
rect 29236 27172 29240 27228
rect 29240 27172 29296 27228
rect 29296 27172 29300 27228
rect 29236 27168 29300 27172
rect 4176 26684 4240 26688
rect 4176 26628 4180 26684
rect 4180 26628 4236 26684
rect 4236 26628 4240 26684
rect 4176 26624 4240 26628
rect 4256 26684 4320 26688
rect 4256 26628 4260 26684
rect 4260 26628 4316 26684
rect 4316 26628 4320 26684
rect 4256 26624 4320 26628
rect 4336 26684 4400 26688
rect 4336 26628 4340 26684
rect 4340 26628 4396 26684
rect 4396 26628 4400 26684
rect 4336 26624 4400 26628
rect 4416 26684 4480 26688
rect 4416 26628 4420 26684
rect 4420 26628 4476 26684
rect 4476 26628 4480 26684
rect 4416 26624 4480 26628
rect 4496 26684 4560 26688
rect 4496 26628 4500 26684
rect 4500 26628 4556 26684
rect 4556 26628 4560 26684
rect 4496 26624 4560 26628
rect 10176 26684 10240 26688
rect 10176 26628 10180 26684
rect 10180 26628 10236 26684
rect 10236 26628 10240 26684
rect 10176 26624 10240 26628
rect 10256 26684 10320 26688
rect 10256 26628 10260 26684
rect 10260 26628 10316 26684
rect 10316 26628 10320 26684
rect 10256 26624 10320 26628
rect 10336 26684 10400 26688
rect 10336 26628 10340 26684
rect 10340 26628 10396 26684
rect 10396 26628 10400 26684
rect 10336 26624 10400 26628
rect 10416 26684 10480 26688
rect 10416 26628 10420 26684
rect 10420 26628 10476 26684
rect 10476 26628 10480 26684
rect 10416 26624 10480 26628
rect 10496 26684 10560 26688
rect 10496 26628 10500 26684
rect 10500 26628 10556 26684
rect 10556 26628 10560 26684
rect 10496 26624 10560 26628
rect 16176 26684 16240 26688
rect 16176 26628 16180 26684
rect 16180 26628 16236 26684
rect 16236 26628 16240 26684
rect 16176 26624 16240 26628
rect 16256 26684 16320 26688
rect 16256 26628 16260 26684
rect 16260 26628 16316 26684
rect 16316 26628 16320 26684
rect 16256 26624 16320 26628
rect 16336 26684 16400 26688
rect 16336 26628 16340 26684
rect 16340 26628 16396 26684
rect 16396 26628 16400 26684
rect 16336 26624 16400 26628
rect 16416 26684 16480 26688
rect 16416 26628 16420 26684
rect 16420 26628 16476 26684
rect 16476 26628 16480 26684
rect 16416 26624 16480 26628
rect 16496 26684 16560 26688
rect 16496 26628 16500 26684
rect 16500 26628 16556 26684
rect 16556 26628 16560 26684
rect 16496 26624 16560 26628
rect 22176 26684 22240 26688
rect 22176 26628 22180 26684
rect 22180 26628 22236 26684
rect 22236 26628 22240 26684
rect 22176 26624 22240 26628
rect 22256 26684 22320 26688
rect 22256 26628 22260 26684
rect 22260 26628 22316 26684
rect 22316 26628 22320 26684
rect 22256 26624 22320 26628
rect 22336 26684 22400 26688
rect 22336 26628 22340 26684
rect 22340 26628 22396 26684
rect 22396 26628 22400 26684
rect 22336 26624 22400 26628
rect 22416 26684 22480 26688
rect 22416 26628 22420 26684
rect 22420 26628 22476 26684
rect 22476 26628 22480 26684
rect 22416 26624 22480 26628
rect 22496 26684 22560 26688
rect 22496 26628 22500 26684
rect 22500 26628 22556 26684
rect 22556 26628 22560 26684
rect 22496 26624 22560 26628
rect 28176 26684 28240 26688
rect 28176 26628 28180 26684
rect 28180 26628 28236 26684
rect 28236 26628 28240 26684
rect 28176 26624 28240 26628
rect 28256 26684 28320 26688
rect 28256 26628 28260 26684
rect 28260 26628 28316 26684
rect 28316 26628 28320 26684
rect 28256 26624 28320 26628
rect 28336 26684 28400 26688
rect 28336 26628 28340 26684
rect 28340 26628 28396 26684
rect 28396 26628 28400 26684
rect 28336 26624 28400 26628
rect 28416 26684 28480 26688
rect 28416 26628 28420 26684
rect 28420 26628 28476 26684
rect 28476 26628 28480 26684
rect 28416 26624 28480 26628
rect 28496 26684 28560 26688
rect 28496 26628 28500 26684
rect 28500 26628 28556 26684
rect 28556 26628 28560 26684
rect 28496 26624 28560 26628
rect 18644 26344 18708 26348
rect 18644 26288 18694 26344
rect 18694 26288 18708 26344
rect 18644 26284 18708 26288
rect 4916 26140 4980 26144
rect 4916 26084 4920 26140
rect 4920 26084 4976 26140
rect 4976 26084 4980 26140
rect 4916 26080 4980 26084
rect 4996 26140 5060 26144
rect 4996 26084 5000 26140
rect 5000 26084 5056 26140
rect 5056 26084 5060 26140
rect 4996 26080 5060 26084
rect 5076 26140 5140 26144
rect 5076 26084 5080 26140
rect 5080 26084 5136 26140
rect 5136 26084 5140 26140
rect 5076 26080 5140 26084
rect 5156 26140 5220 26144
rect 5156 26084 5160 26140
rect 5160 26084 5216 26140
rect 5216 26084 5220 26140
rect 5156 26080 5220 26084
rect 5236 26140 5300 26144
rect 5236 26084 5240 26140
rect 5240 26084 5296 26140
rect 5296 26084 5300 26140
rect 5236 26080 5300 26084
rect 10916 26140 10980 26144
rect 10916 26084 10920 26140
rect 10920 26084 10976 26140
rect 10976 26084 10980 26140
rect 10916 26080 10980 26084
rect 10996 26140 11060 26144
rect 10996 26084 11000 26140
rect 11000 26084 11056 26140
rect 11056 26084 11060 26140
rect 10996 26080 11060 26084
rect 11076 26140 11140 26144
rect 11076 26084 11080 26140
rect 11080 26084 11136 26140
rect 11136 26084 11140 26140
rect 11076 26080 11140 26084
rect 11156 26140 11220 26144
rect 11156 26084 11160 26140
rect 11160 26084 11216 26140
rect 11216 26084 11220 26140
rect 11156 26080 11220 26084
rect 11236 26140 11300 26144
rect 11236 26084 11240 26140
rect 11240 26084 11296 26140
rect 11296 26084 11300 26140
rect 11236 26080 11300 26084
rect 16916 26140 16980 26144
rect 16916 26084 16920 26140
rect 16920 26084 16976 26140
rect 16976 26084 16980 26140
rect 16916 26080 16980 26084
rect 16996 26140 17060 26144
rect 16996 26084 17000 26140
rect 17000 26084 17056 26140
rect 17056 26084 17060 26140
rect 16996 26080 17060 26084
rect 17076 26140 17140 26144
rect 17076 26084 17080 26140
rect 17080 26084 17136 26140
rect 17136 26084 17140 26140
rect 17076 26080 17140 26084
rect 17156 26140 17220 26144
rect 17156 26084 17160 26140
rect 17160 26084 17216 26140
rect 17216 26084 17220 26140
rect 17156 26080 17220 26084
rect 17236 26140 17300 26144
rect 17236 26084 17240 26140
rect 17240 26084 17296 26140
rect 17296 26084 17300 26140
rect 17236 26080 17300 26084
rect 22916 26140 22980 26144
rect 22916 26084 22920 26140
rect 22920 26084 22976 26140
rect 22976 26084 22980 26140
rect 22916 26080 22980 26084
rect 22996 26140 23060 26144
rect 22996 26084 23000 26140
rect 23000 26084 23056 26140
rect 23056 26084 23060 26140
rect 22996 26080 23060 26084
rect 23076 26140 23140 26144
rect 23076 26084 23080 26140
rect 23080 26084 23136 26140
rect 23136 26084 23140 26140
rect 23076 26080 23140 26084
rect 23156 26140 23220 26144
rect 23156 26084 23160 26140
rect 23160 26084 23216 26140
rect 23216 26084 23220 26140
rect 23156 26080 23220 26084
rect 23236 26140 23300 26144
rect 23236 26084 23240 26140
rect 23240 26084 23296 26140
rect 23296 26084 23300 26140
rect 23236 26080 23300 26084
rect 28916 26140 28980 26144
rect 28916 26084 28920 26140
rect 28920 26084 28976 26140
rect 28976 26084 28980 26140
rect 28916 26080 28980 26084
rect 28996 26140 29060 26144
rect 28996 26084 29000 26140
rect 29000 26084 29056 26140
rect 29056 26084 29060 26140
rect 28996 26080 29060 26084
rect 29076 26140 29140 26144
rect 29076 26084 29080 26140
rect 29080 26084 29136 26140
rect 29136 26084 29140 26140
rect 29076 26080 29140 26084
rect 29156 26140 29220 26144
rect 29156 26084 29160 26140
rect 29160 26084 29216 26140
rect 29216 26084 29220 26140
rect 29156 26080 29220 26084
rect 29236 26140 29300 26144
rect 29236 26084 29240 26140
rect 29240 26084 29296 26140
rect 29296 26084 29300 26140
rect 29236 26080 29300 26084
rect 4176 25596 4240 25600
rect 4176 25540 4180 25596
rect 4180 25540 4236 25596
rect 4236 25540 4240 25596
rect 4176 25536 4240 25540
rect 4256 25596 4320 25600
rect 4256 25540 4260 25596
rect 4260 25540 4316 25596
rect 4316 25540 4320 25596
rect 4256 25536 4320 25540
rect 4336 25596 4400 25600
rect 4336 25540 4340 25596
rect 4340 25540 4396 25596
rect 4396 25540 4400 25596
rect 4336 25536 4400 25540
rect 4416 25596 4480 25600
rect 4416 25540 4420 25596
rect 4420 25540 4476 25596
rect 4476 25540 4480 25596
rect 4416 25536 4480 25540
rect 4496 25596 4560 25600
rect 4496 25540 4500 25596
rect 4500 25540 4556 25596
rect 4556 25540 4560 25596
rect 4496 25536 4560 25540
rect 10176 25596 10240 25600
rect 10176 25540 10180 25596
rect 10180 25540 10236 25596
rect 10236 25540 10240 25596
rect 10176 25536 10240 25540
rect 10256 25596 10320 25600
rect 10256 25540 10260 25596
rect 10260 25540 10316 25596
rect 10316 25540 10320 25596
rect 10256 25536 10320 25540
rect 10336 25596 10400 25600
rect 10336 25540 10340 25596
rect 10340 25540 10396 25596
rect 10396 25540 10400 25596
rect 10336 25536 10400 25540
rect 10416 25596 10480 25600
rect 10416 25540 10420 25596
rect 10420 25540 10476 25596
rect 10476 25540 10480 25596
rect 10416 25536 10480 25540
rect 10496 25596 10560 25600
rect 10496 25540 10500 25596
rect 10500 25540 10556 25596
rect 10556 25540 10560 25596
rect 10496 25536 10560 25540
rect 16176 25596 16240 25600
rect 16176 25540 16180 25596
rect 16180 25540 16236 25596
rect 16236 25540 16240 25596
rect 16176 25536 16240 25540
rect 16256 25596 16320 25600
rect 16256 25540 16260 25596
rect 16260 25540 16316 25596
rect 16316 25540 16320 25596
rect 16256 25536 16320 25540
rect 16336 25596 16400 25600
rect 16336 25540 16340 25596
rect 16340 25540 16396 25596
rect 16396 25540 16400 25596
rect 16336 25536 16400 25540
rect 16416 25596 16480 25600
rect 16416 25540 16420 25596
rect 16420 25540 16476 25596
rect 16476 25540 16480 25596
rect 16416 25536 16480 25540
rect 16496 25596 16560 25600
rect 16496 25540 16500 25596
rect 16500 25540 16556 25596
rect 16556 25540 16560 25596
rect 16496 25536 16560 25540
rect 22176 25596 22240 25600
rect 22176 25540 22180 25596
rect 22180 25540 22236 25596
rect 22236 25540 22240 25596
rect 22176 25536 22240 25540
rect 22256 25596 22320 25600
rect 22256 25540 22260 25596
rect 22260 25540 22316 25596
rect 22316 25540 22320 25596
rect 22256 25536 22320 25540
rect 22336 25596 22400 25600
rect 22336 25540 22340 25596
rect 22340 25540 22396 25596
rect 22396 25540 22400 25596
rect 22336 25536 22400 25540
rect 22416 25596 22480 25600
rect 22416 25540 22420 25596
rect 22420 25540 22476 25596
rect 22476 25540 22480 25596
rect 22416 25536 22480 25540
rect 22496 25596 22560 25600
rect 22496 25540 22500 25596
rect 22500 25540 22556 25596
rect 22556 25540 22560 25596
rect 22496 25536 22560 25540
rect 28176 25596 28240 25600
rect 28176 25540 28180 25596
rect 28180 25540 28236 25596
rect 28236 25540 28240 25596
rect 28176 25536 28240 25540
rect 28256 25596 28320 25600
rect 28256 25540 28260 25596
rect 28260 25540 28316 25596
rect 28316 25540 28320 25596
rect 28256 25536 28320 25540
rect 28336 25596 28400 25600
rect 28336 25540 28340 25596
rect 28340 25540 28396 25596
rect 28396 25540 28400 25596
rect 28336 25536 28400 25540
rect 28416 25596 28480 25600
rect 28416 25540 28420 25596
rect 28420 25540 28476 25596
rect 28476 25540 28480 25596
rect 28416 25536 28480 25540
rect 28496 25596 28560 25600
rect 28496 25540 28500 25596
rect 28500 25540 28556 25596
rect 28556 25540 28560 25596
rect 28496 25536 28560 25540
rect 4916 25052 4980 25056
rect 4916 24996 4920 25052
rect 4920 24996 4976 25052
rect 4976 24996 4980 25052
rect 4916 24992 4980 24996
rect 4996 25052 5060 25056
rect 4996 24996 5000 25052
rect 5000 24996 5056 25052
rect 5056 24996 5060 25052
rect 4996 24992 5060 24996
rect 5076 25052 5140 25056
rect 5076 24996 5080 25052
rect 5080 24996 5136 25052
rect 5136 24996 5140 25052
rect 5076 24992 5140 24996
rect 5156 25052 5220 25056
rect 5156 24996 5160 25052
rect 5160 24996 5216 25052
rect 5216 24996 5220 25052
rect 5156 24992 5220 24996
rect 5236 25052 5300 25056
rect 5236 24996 5240 25052
rect 5240 24996 5296 25052
rect 5296 24996 5300 25052
rect 5236 24992 5300 24996
rect 10916 25052 10980 25056
rect 10916 24996 10920 25052
rect 10920 24996 10976 25052
rect 10976 24996 10980 25052
rect 10916 24992 10980 24996
rect 10996 25052 11060 25056
rect 10996 24996 11000 25052
rect 11000 24996 11056 25052
rect 11056 24996 11060 25052
rect 10996 24992 11060 24996
rect 11076 25052 11140 25056
rect 11076 24996 11080 25052
rect 11080 24996 11136 25052
rect 11136 24996 11140 25052
rect 11076 24992 11140 24996
rect 11156 25052 11220 25056
rect 11156 24996 11160 25052
rect 11160 24996 11216 25052
rect 11216 24996 11220 25052
rect 11156 24992 11220 24996
rect 11236 25052 11300 25056
rect 11236 24996 11240 25052
rect 11240 24996 11296 25052
rect 11296 24996 11300 25052
rect 11236 24992 11300 24996
rect 16916 25052 16980 25056
rect 16916 24996 16920 25052
rect 16920 24996 16976 25052
rect 16976 24996 16980 25052
rect 16916 24992 16980 24996
rect 16996 25052 17060 25056
rect 16996 24996 17000 25052
rect 17000 24996 17056 25052
rect 17056 24996 17060 25052
rect 16996 24992 17060 24996
rect 17076 25052 17140 25056
rect 17076 24996 17080 25052
rect 17080 24996 17136 25052
rect 17136 24996 17140 25052
rect 17076 24992 17140 24996
rect 17156 25052 17220 25056
rect 17156 24996 17160 25052
rect 17160 24996 17216 25052
rect 17216 24996 17220 25052
rect 17156 24992 17220 24996
rect 17236 25052 17300 25056
rect 17236 24996 17240 25052
rect 17240 24996 17296 25052
rect 17296 24996 17300 25052
rect 17236 24992 17300 24996
rect 22916 25052 22980 25056
rect 22916 24996 22920 25052
rect 22920 24996 22976 25052
rect 22976 24996 22980 25052
rect 22916 24992 22980 24996
rect 22996 25052 23060 25056
rect 22996 24996 23000 25052
rect 23000 24996 23056 25052
rect 23056 24996 23060 25052
rect 22996 24992 23060 24996
rect 23076 25052 23140 25056
rect 23076 24996 23080 25052
rect 23080 24996 23136 25052
rect 23136 24996 23140 25052
rect 23076 24992 23140 24996
rect 23156 25052 23220 25056
rect 23156 24996 23160 25052
rect 23160 24996 23216 25052
rect 23216 24996 23220 25052
rect 23156 24992 23220 24996
rect 23236 25052 23300 25056
rect 23236 24996 23240 25052
rect 23240 24996 23296 25052
rect 23296 24996 23300 25052
rect 23236 24992 23300 24996
rect 28916 25052 28980 25056
rect 28916 24996 28920 25052
rect 28920 24996 28976 25052
rect 28976 24996 28980 25052
rect 28916 24992 28980 24996
rect 28996 25052 29060 25056
rect 28996 24996 29000 25052
rect 29000 24996 29056 25052
rect 29056 24996 29060 25052
rect 28996 24992 29060 24996
rect 29076 25052 29140 25056
rect 29076 24996 29080 25052
rect 29080 24996 29136 25052
rect 29136 24996 29140 25052
rect 29076 24992 29140 24996
rect 29156 25052 29220 25056
rect 29156 24996 29160 25052
rect 29160 24996 29216 25052
rect 29216 24996 29220 25052
rect 29156 24992 29220 24996
rect 29236 25052 29300 25056
rect 29236 24996 29240 25052
rect 29240 24996 29296 25052
rect 29296 24996 29300 25052
rect 29236 24992 29300 24996
rect 4176 24508 4240 24512
rect 4176 24452 4180 24508
rect 4180 24452 4236 24508
rect 4236 24452 4240 24508
rect 4176 24448 4240 24452
rect 4256 24508 4320 24512
rect 4256 24452 4260 24508
rect 4260 24452 4316 24508
rect 4316 24452 4320 24508
rect 4256 24448 4320 24452
rect 4336 24508 4400 24512
rect 4336 24452 4340 24508
rect 4340 24452 4396 24508
rect 4396 24452 4400 24508
rect 4336 24448 4400 24452
rect 4416 24508 4480 24512
rect 4416 24452 4420 24508
rect 4420 24452 4476 24508
rect 4476 24452 4480 24508
rect 4416 24448 4480 24452
rect 4496 24508 4560 24512
rect 4496 24452 4500 24508
rect 4500 24452 4556 24508
rect 4556 24452 4560 24508
rect 4496 24448 4560 24452
rect 10176 24508 10240 24512
rect 10176 24452 10180 24508
rect 10180 24452 10236 24508
rect 10236 24452 10240 24508
rect 10176 24448 10240 24452
rect 10256 24508 10320 24512
rect 10256 24452 10260 24508
rect 10260 24452 10316 24508
rect 10316 24452 10320 24508
rect 10256 24448 10320 24452
rect 10336 24508 10400 24512
rect 10336 24452 10340 24508
rect 10340 24452 10396 24508
rect 10396 24452 10400 24508
rect 10336 24448 10400 24452
rect 10416 24508 10480 24512
rect 10416 24452 10420 24508
rect 10420 24452 10476 24508
rect 10476 24452 10480 24508
rect 10416 24448 10480 24452
rect 10496 24508 10560 24512
rect 10496 24452 10500 24508
rect 10500 24452 10556 24508
rect 10556 24452 10560 24508
rect 10496 24448 10560 24452
rect 16176 24508 16240 24512
rect 16176 24452 16180 24508
rect 16180 24452 16236 24508
rect 16236 24452 16240 24508
rect 16176 24448 16240 24452
rect 16256 24508 16320 24512
rect 16256 24452 16260 24508
rect 16260 24452 16316 24508
rect 16316 24452 16320 24508
rect 16256 24448 16320 24452
rect 16336 24508 16400 24512
rect 16336 24452 16340 24508
rect 16340 24452 16396 24508
rect 16396 24452 16400 24508
rect 16336 24448 16400 24452
rect 16416 24508 16480 24512
rect 16416 24452 16420 24508
rect 16420 24452 16476 24508
rect 16476 24452 16480 24508
rect 16416 24448 16480 24452
rect 16496 24508 16560 24512
rect 16496 24452 16500 24508
rect 16500 24452 16556 24508
rect 16556 24452 16560 24508
rect 16496 24448 16560 24452
rect 22176 24508 22240 24512
rect 22176 24452 22180 24508
rect 22180 24452 22236 24508
rect 22236 24452 22240 24508
rect 22176 24448 22240 24452
rect 22256 24508 22320 24512
rect 22256 24452 22260 24508
rect 22260 24452 22316 24508
rect 22316 24452 22320 24508
rect 22256 24448 22320 24452
rect 22336 24508 22400 24512
rect 22336 24452 22340 24508
rect 22340 24452 22396 24508
rect 22396 24452 22400 24508
rect 22336 24448 22400 24452
rect 22416 24508 22480 24512
rect 22416 24452 22420 24508
rect 22420 24452 22476 24508
rect 22476 24452 22480 24508
rect 22416 24448 22480 24452
rect 22496 24508 22560 24512
rect 22496 24452 22500 24508
rect 22500 24452 22556 24508
rect 22556 24452 22560 24508
rect 22496 24448 22560 24452
rect 28176 24508 28240 24512
rect 28176 24452 28180 24508
rect 28180 24452 28236 24508
rect 28236 24452 28240 24508
rect 28176 24448 28240 24452
rect 28256 24508 28320 24512
rect 28256 24452 28260 24508
rect 28260 24452 28316 24508
rect 28316 24452 28320 24508
rect 28256 24448 28320 24452
rect 28336 24508 28400 24512
rect 28336 24452 28340 24508
rect 28340 24452 28396 24508
rect 28396 24452 28400 24508
rect 28336 24448 28400 24452
rect 28416 24508 28480 24512
rect 28416 24452 28420 24508
rect 28420 24452 28476 24508
rect 28476 24452 28480 24508
rect 28416 24448 28480 24452
rect 28496 24508 28560 24512
rect 28496 24452 28500 24508
rect 28500 24452 28556 24508
rect 28556 24452 28560 24508
rect 28496 24448 28560 24452
rect 4916 23964 4980 23968
rect 4916 23908 4920 23964
rect 4920 23908 4976 23964
rect 4976 23908 4980 23964
rect 4916 23904 4980 23908
rect 4996 23964 5060 23968
rect 4996 23908 5000 23964
rect 5000 23908 5056 23964
rect 5056 23908 5060 23964
rect 4996 23904 5060 23908
rect 5076 23964 5140 23968
rect 5076 23908 5080 23964
rect 5080 23908 5136 23964
rect 5136 23908 5140 23964
rect 5076 23904 5140 23908
rect 5156 23964 5220 23968
rect 5156 23908 5160 23964
rect 5160 23908 5216 23964
rect 5216 23908 5220 23964
rect 5156 23904 5220 23908
rect 5236 23964 5300 23968
rect 5236 23908 5240 23964
rect 5240 23908 5296 23964
rect 5296 23908 5300 23964
rect 5236 23904 5300 23908
rect 10916 23964 10980 23968
rect 10916 23908 10920 23964
rect 10920 23908 10976 23964
rect 10976 23908 10980 23964
rect 10916 23904 10980 23908
rect 10996 23964 11060 23968
rect 10996 23908 11000 23964
rect 11000 23908 11056 23964
rect 11056 23908 11060 23964
rect 10996 23904 11060 23908
rect 11076 23964 11140 23968
rect 11076 23908 11080 23964
rect 11080 23908 11136 23964
rect 11136 23908 11140 23964
rect 11076 23904 11140 23908
rect 11156 23964 11220 23968
rect 11156 23908 11160 23964
rect 11160 23908 11216 23964
rect 11216 23908 11220 23964
rect 11156 23904 11220 23908
rect 11236 23964 11300 23968
rect 11236 23908 11240 23964
rect 11240 23908 11296 23964
rect 11296 23908 11300 23964
rect 11236 23904 11300 23908
rect 16916 23964 16980 23968
rect 16916 23908 16920 23964
rect 16920 23908 16976 23964
rect 16976 23908 16980 23964
rect 16916 23904 16980 23908
rect 16996 23964 17060 23968
rect 16996 23908 17000 23964
rect 17000 23908 17056 23964
rect 17056 23908 17060 23964
rect 16996 23904 17060 23908
rect 17076 23964 17140 23968
rect 17076 23908 17080 23964
rect 17080 23908 17136 23964
rect 17136 23908 17140 23964
rect 17076 23904 17140 23908
rect 17156 23964 17220 23968
rect 17156 23908 17160 23964
rect 17160 23908 17216 23964
rect 17216 23908 17220 23964
rect 17156 23904 17220 23908
rect 17236 23964 17300 23968
rect 17236 23908 17240 23964
rect 17240 23908 17296 23964
rect 17296 23908 17300 23964
rect 17236 23904 17300 23908
rect 22916 23964 22980 23968
rect 22916 23908 22920 23964
rect 22920 23908 22976 23964
rect 22976 23908 22980 23964
rect 22916 23904 22980 23908
rect 22996 23964 23060 23968
rect 22996 23908 23000 23964
rect 23000 23908 23056 23964
rect 23056 23908 23060 23964
rect 22996 23904 23060 23908
rect 23076 23964 23140 23968
rect 23076 23908 23080 23964
rect 23080 23908 23136 23964
rect 23136 23908 23140 23964
rect 23076 23904 23140 23908
rect 23156 23964 23220 23968
rect 23156 23908 23160 23964
rect 23160 23908 23216 23964
rect 23216 23908 23220 23964
rect 23156 23904 23220 23908
rect 23236 23964 23300 23968
rect 23236 23908 23240 23964
rect 23240 23908 23296 23964
rect 23296 23908 23300 23964
rect 23236 23904 23300 23908
rect 28916 23964 28980 23968
rect 28916 23908 28920 23964
rect 28920 23908 28976 23964
rect 28976 23908 28980 23964
rect 28916 23904 28980 23908
rect 28996 23964 29060 23968
rect 28996 23908 29000 23964
rect 29000 23908 29056 23964
rect 29056 23908 29060 23964
rect 28996 23904 29060 23908
rect 29076 23964 29140 23968
rect 29076 23908 29080 23964
rect 29080 23908 29136 23964
rect 29136 23908 29140 23964
rect 29076 23904 29140 23908
rect 29156 23964 29220 23968
rect 29156 23908 29160 23964
rect 29160 23908 29216 23964
rect 29216 23908 29220 23964
rect 29156 23904 29220 23908
rect 29236 23964 29300 23968
rect 29236 23908 29240 23964
rect 29240 23908 29296 23964
rect 29296 23908 29300 23964
rect 29236 23904 29300 23908
rect 15332 23564 15396 23628
rect 4176 23420 4240 23424
rect 4176 23364 4180 23420
rect 4180 23364 4236 23420
rect 4236 23364 4240 23420
rect 4176 23360 4240 23364
rect 4256 23420 4320 23424
rect 4256 23364 4260 23420
rect 4260 23364 4316 23420
rect 4316 23364 4320 23420
rect 4256 23360 4320 23364
rect 4336 23420 4400 23424
rect 4336 23364 4340 23420
rect 4340 23364 4396 23420
rect 4396 23364 4400 23420
rect 4336 23360 4400 23364
rect 4416 23420 4480 23424
rect 4416 23364 4420 23420
rect 4420 23364 4476 23420
rect 4476 23364 4480 23420
rect 4416 23360 4480 23364
rect 4496 23420 4560 23424
rect 4496 23364 4500 23420
rect 4500 23364 4556 23420
rect 4556 23364 4560 23420
rect 4496 23360 4560 23364
rect 10176 23420 10240 23424
rect 10176 23364 10180 23420
rect 10180 23364 10236 23420
rect 10236 23364 10240 23420
rect 10176 23360 10240 23364
rect 10256 23420 10320 23424
rect 10256 23364 10260 23420
rect 10260 23364 10316 23420
rect 10316 23364 10320 23420
rect 10256 23360 10320 23364
rect 10336 23420 10400 23424
rect 10336 23364 10340 23420
rect 10340 23364 10396 23420
rect 10396 23364 10400 23420
rect 10336 23360 10400 23364
rect 10416 23420 10480 23424
rect 10416 23364 10420 23420
rect 10420 23364 10476 23420
rect 10476 23364 10480 23420
rect 10416 23360 10480 23364
rect 10496 23420 10560 23424
rect 10496 23364 10500 23420
rect 10500 23364 10556 23420
rect 10556 23364 10560 23420
rect 10496 23360 10560 23364
rect 16176 23420 16240 23424
rect 16176 23364 16180 23420
rect 16180 23364 16236 23420
rect 16236 23364 16240 23420
rect 16176 23360 16240 23364
rect 16256 23420 16320 23424
rect 16256 23364 16260 23420
rect 16260 23364 16316 23420
rect 16316 23364 16320 23420
rect 16256 23360 16320 23364
rect 16336 23420 16400 23424
rect 16336 23364 16340 23420
rect 16340 23364 16396 23420
rect 16396 23364 16400 23420
rect 16336 23360 16400 23364
rect 16416 23420 16480 23424
rect 16416 23364 16420 23420
rect 16420 23364 16476 23420
rect 16476 23364 16480 23420
rect 16416 23360 16480 23364
rect 16496 23420 16560 23424
rect 16496 23364 16500 23420
rect 16500 23364 16556 23420
rect 16556 23364 16560 23420
rect 16496 23360 16560 23364
rect 22176 23420 22240 23424
rect 22176 23364 22180 23420
rect 22180 23364 22236 23420
rect 22236 23364 22240 23420
rect 22176 23360 22240 23364
rect 22256 23420 22320 23424
rect 22256 23364 22260 23420
rect 22260 23364 22316 23420
rect 22316 23364 22320 23420
rect 22256 23360 22320 23364
rect 22336 23420 22400 23424
rect 22336 23364 22340 23420
rect 22340 23364 22396 23420
rect 22396 23364 22400 23420
rect 22336 23360 22400 23364
rect 22416 23420 22480 23424
rect 22416 23364 22420 23420
rect 22420 23364 22476 23420
rect 22476 23364 22480 23420
rect 22416 23360 22480 23364
rect 22496 23420 22560 23424
rect 22496 23364 22500 23420
rect 22500 23364 22556 23420
rect 22556 23364 22560 23420
rect 22496 23360 22560 23364
rect 28176 23420 28240 23424
rect 28176 23364 28180 23420
rect 28180 23364 28236 23420
rect 28236 23364 28240 23420
rect 28176 23360 28240 23364
rect 28256 23420 28320 23424
rect 28256 23364 28260 23420
rect 28260 23364 28316 23420
rect 28316 23364 28320 23420
rect 28256 23360 28320 23364
rect 28336 23420 28400 23424
rect 28336 23364 28340 23420
rect 28340 23364 28396 23420
rect 28396 23364 28400 23420
rect 28336 23360 28400 23364
rect 28416 23420 28480 23424
rect 28416 23364 28420 23420
rect 28420 23364 28476 23420
rect 28476 23364 28480 23420
rect 28416 23360 28480 23364
rect 28496 23420 28560 23424
rect 28496 23364 28500 23420
rect 28500 23364 28556 23420
rect 28556 23364 28560 23420
rect 28496 23360 28560 23364
rect 4916 22876 4980 22880
rect 4916 22820 4920 22876
rect 4920 22820 4976 22876
rect 4976 22820 4980 22876
rect 4916 22816 4980 22820
rect 4996 22876 5060 22880
rect 4996 22820 5000 22876
rect 5000 22820 5056 22876
rect 5056 22820 5060 22876
rect 4996 22816 5060 22820
rect 5076 22876 5140 22880
rect 5076 22820 5080 22876
rect 5080 22820 5136 22876
rect 5136 22820 5140 22876
rect 5076 22816 5140 22820
rect 5156 22876 5220 22880
rect 5156 22820 5160 22876
rect 5160 22820 5216 22876
rect 5216 22820 5220 22876
rect 5156 22816 5220 22820
rect 5236 22876 5300 22880
rect 5236 22820 5240 22876
rect 5240 22820 5296 22876
rect 5296 22820 5300 22876
rect 5236 22816 5300 22820
rect 10916 22876 10980 22880
rect 10916 22820 10920 22876
rect 10920 22820 10976 22876
rect 10976 22820 10980 22876
rect 10916 22816 10980 22820
rect 10996 22876 11060 22880
rect 10996 22820 11000 22876
rect 11000 22820 11056 22876
rect 11056 22820 11060 22876
rect 10996 22816 11060 22820
rect 11076 22876 11140 22880
rect 11076 22820 11080 22876
rect 11080 22820 11136 22876
rect 11136 22820 11140 22876
rect 11076 22816 11140 22820
rect 11156 22876 11220 22880
rect 11156 22820 11160 22876
rect 11160 22820 11216 22876
rect 11216 22820 11220 22876
rect 11156 22816 11220 22820
rect 11236 22876 11300 22880
rect 11236 22820 11240 22876
rect 11240 22820 11296 22876
rect 11296 22820 11300 22876
rect 11236 22816 11300 22820
rect 16916 22876 16980 22880
rect 16916 22820 16920 22876
rect 16920 22820 16976 22876
rect 16976 22820 16980 22876
rect 16916 22816 16980 22820
rect 16996 22876 17060 22880
rect 16996 22820 17000 22876
rect 17000 22820 17056 22876
rect 17056 22820 17060 22876
rect 16996 22816 17060 22820
rect 17076 22876 17140 22880
rect 17076 22820 17080 22876
rect 17080 22820 17136 22876
rect 17136 22820 17140 22876
rect 17076 22816 17140 22820
rect 17156 22876 17220 22880
rect 17156 22820 17160 22876
rect 17160 22820 17216 22876
rect 17216 22820 17220 22876
rect 17156 22816 17220 22820
rect 17236 22876 17300 22880
rect 17236 22820 17240 22876
rect 17240 22820 17296 22876
rect 17296 22820 17300 22876
rect 17236 22816 17300 22820
rect 22916 22876 22980 22880
rect 22916 22820 22920 22876
rect 22920 22820 22976 22876
rect 22976 22820 22980 22876
rect 22916 22816 22980 22820
rect 22996 22876 23060 22880
rect 22996 22820 23000 22876
rect 23000 22820 23056 22876
rect 23056 22820 23060 22876
rect 22996 22816 23060 22820
rect 23076 22876 23140 22880
rect 23076 22820 23080 22876
rect 23080 22820 23136 22876
rect 23136 22820 23140 22876
rect 23076 22816 23140 22820
rect 23156 22876 23220 22880
rect 23156 22820 23160 22876
rect 23160 22820 23216 22876
rect 23216 22820 23220 22876
rect 23156 22816 23220 22820
rect 23236 22876 23300 22880
rect 23236 22820 23240 22876
rect 23240 22820 23296 22876
rect 23296 22820 23300 22876
rect 23236 22816 23300 22820
rect 28916 22876 28980 22880
rect 28916 22820 28920 22876
rect 28920 22820 28976 22876
rect 28976 22820 28980 22876
rect 28916 22816 28980 22820
rect 28996 22876 29060 22880
rect 28996 22820 29000 22876
rect 29000 22820 29056 22876
rect 29056 22820 29060 22876
rect 28996 22816 29060 22820
rect 29076 22876 29140 22880
rect 29076 22820 29080 22876
rect 29080 22820 29136 22876
rect 29136 22820 29140 22876
rect 29076 22816 29140 22820
rect 29156 22876 29220 22880
rect 29156 22820 29160 22876
rect 29160 22820 29216 22876
rect 29216 22820 29220 22876
rect 29156 22816 29220 22820
rect 29236 22876 29300 22880
rect 29236 22820 29240 22876
rect 29240 22820 29296 22876
rect 29296 22820 29300 22876
rect 29236 22816 29300 22820
rect 4176 22332 4240 22336
rect 4176 22276 4180 22332
rect 4180 22276 4236 22332
rect 4236 22276 4240 22332
rect 4176 22272 4240 22276
rect 4256 22332 4320 22336
rect 4256 22276 4260 22332
rect 4260 22276 4316 22332
rect 4316 22276 4320 22332
rect 4256 22272 4320 22276
rect 4336 22332 4400 22336
rect 4336 22276 4340 22332
rect 4340 22276 4396 22332
rect 4396 22276 4400 22332
rect 4336 22272 4400 22276
rect 4416 22332 4480 22336
rect 4416 22276 4420 22332
rect 4420 22276 4476 22332
rect 4476 22276 4480 22332
rect 4416 22272 4480 22276
rect 4496 22332 4560 22336
rect 4496 22276 4500 22332
rect 4500 22276 4556 22332
rect 4556 22276 4560 22332
rect 4496 22272 4560 22276
rect 10176 22332 10240 22336
rect 10176 22276 10180 22332
rect 10180 22276 10236 22332
rect 10236 22276 10240 22332
rect 10176 22272 10240 22276
rect 10256 22332 10320 22336
rect 10256 22276 10260 22332
rect 10260 22276 10316 22332
rect 10316 22276 10320 22332
rect 10256 22272 10320 22276
rect 10336 22332 10400 22336
rect 10336 22276 10340 22332
rect 10340 22276 10396 22332
rect 10396 22276 10400 22332
rect 10336 22272 10400 22276
rect 10416 22332 10480 22336
rect 10416 22276 10420 22332
rect 10420 22276 10476 22332
rect 10476 22276 10480 22332
rect 10416 22272 10480 22276
rect 10496 22332 10560 22336
rect 10496 22276 10500 22332
rect 10500 22276 10556 22332
rect 10556 22276 10560 22332
rect 10496 22272 10560 22276
rect 16176 22332 16240 22336
rect 16176 22276 16180 22332
rect 16180 22276 16236 22332
rect 16236 22276 16240 22332
rect 16176 22272 16240 22276
rect 16256 22332 16320 22336
rect 16256 22276 16260 22332
rect 16260 22276 16316 22332
rect 16316 22276 16320 22332
rect 16256 22272 16320 22276
rect 16336 22332 16400 22336
rect 16336 22276 16340 22332
rect 16340 22276 16396 22332
rect 16396 22276 16400 22332
rect 16336 22272 16400 22276
rect 16416 22332 16480 22336
rect 16416 22276 16420 22332
rect 16420 22276 16476 22332
rect 16476 22276 16480 22332
rect 16416 22272 16480 22276
rect 16496 22332 16560 22336
rect 16496 22276 16500 22332
rect 16500 22276 16556 22332
rect 16556 22276 16560 22332
rect 16496 22272 16560 22276
rect 22176 22332 22240 22336
rect 22176 22276 22180 22332
rect 22180 22276 22236 22332
rect 22236 22276 22240 22332
rect 22176 22272 22240 22276
rect 22256 22332 22320 22336
rect 22256 22276 22260 22332
rect 22260 22276 22316 22332
rect 22316 22276 22320 22332
rect 22256 22272 22320 22276
rect 22336 22332 22400 22336
rect 22336 22276 22340 22332
rect 22340 22276 22396 22332
rect 22396 22276 22400 22332
rect 22336 22272 22400 22276
rect 22416 22332 22480 22336
rect 22416 22276 22420 22332
rect 22420 22276 22476 22332
rect 22476 22276 22480 22332
rect 22416 22272 22480 22276
rect 22496 22332 22560 22336
rect 22496 22276 22500 22332
rect 22500 22276 22556 22332
rect 22556 22276 22560 22332
rect 22496 22272 22560 22276
rect 28176 22332 28240 22336
rect 28176 22276 28180 22332
rect 28180 22276 28236 22332
rect 28236 22276 28240 22332
rect 28176 22272 28240 22276
rect 28256 22332 28320 22336
rect 28256 22276 28260 22332
rect 28260 22276 28316 22332
rect 28316 22276 28320 22332
rect 28256 22272 28320 22276
rect 28336 22332 28400 22336
rect 28336 22276 28340 22332
rect 28340 22276 28396 22332
rect 28396 22276 28400 22332
rect 28336 22272 28400 22276
rect 28416 22332 28480 22336
rect 28416 22276 28420 22332
rect 28420 22276 28476 22332
rect 28476 22276 28480 22332
rect 28416 22272 28480 22276
rect 28496 22332 28560 22336
rect 28496 22276 28500 22332
rect 28500 22276 28556 22332
rect 28556 22276 28560 22332
rect 28496 22272 28560 22276
rect 24348 21932 24412 21996
rect 4916 21788 4980 21792
rect 4916 21732 4920 21788
rect 4920 21732 4976 21788
rect 4976 21732 4980 21788
rect 4916 21728 4980 21732
rect 4996 21788 5060 21792
rect 4996 21732 5000 21788
rect 5000 21732 5056 21788
rect 5056 21732 5060 21788
rect 4996 21728 5060 21732
rect 5076 21788 5140 21792
rect 5076 21732 5080 21788
rect 5080 21732 5136 21788
rect 5136 21732 5140 21788
rect 5076 21728 5140 21732
rect 5156 21788 5220 21792
rect 5156 21732 5160 21788
rect 5160 21732 5216 21788
rect 5216 21732 5220 21788
rect 5156 21728 5220 21732
rect 5236 21788 5300 21792
rect 5236 21732 5240 21788
rect 5240 21732 5296 21788
rect 5296 21732 5300 21788
rect 5236 21728 5300 21732
rect 10916 21788 10980 21792
rect 10916 21732 10920 21788
rect 10920 21732 10976 21788
rect 10976 21732 10980 21788
rect 10916 21728 10980 21732
rect 10996 21788 11060 21792
rect 10996 21732 11000 21788
rect 11000 21732 11056 21788
rect 11056 21732 11060 21788
rect 10996 21728 11060 21732
rect 11076 21788 11140 21792
rect 11076 21732 11080 21788
rect 11080 21732 11136 21788
rect 11136 21732 11140 21788
rect 11076 21728 11140 21732
rect 11156 21788 11220 21792
rect 11156 21732 11160 21788
rect 11160 21732 11216 21788
rect 11216 21732 11220 21788
rect 11156 21728 11220 21732
rect 11236 21788 11300 21792
rect 11236 21732 11240 21788
rect 11240 21732 11296 21788
rect 11296 21732 11300 21788
rect 11236 21728 11300 21732
rect 16916 21788 16980 21792
rect 16916 21732 16920 21788
rect 16920 21732 16976 21788
rect 16976 21732 16980 21788
rect 16916 21728 16980 21732
rect 16996 21788 17060 21792
rect 16996 21732 17000 21788
rect 17000 21732 17056 21788
rect 17056 21732 17060 21788
rect 16996 21728 17060 21732
rect 17076 21788 17140 21792
rect 17076 21732 17080 21788
rect 17080 21732 17136 21788
rect 17136 21732 17140 21788
rect 17076 21728 17140 21732
rect 17156 21788 17220 21792
rect 17156 21732 17160 21788
rect 17160 21732 17216 21788
rect 17216 21732 17220 21788
rect 17156 21728 17220 21732
rect 17236 21788 17300 21792
rect 17236 21732 17240 21788
rect 17240 21732 17296 21788
rect 17296 21732 17300 21788
rect 17236 21728 17300 21732
rect 22916 21788 22980 21792
rect 22916 21732 22920 21788
rect 22920 21732 22976 21788
rect 22976 21732 22980 21788
rect 22916 21728 22980 21732
rect 22996 21788 23060 21792
rect 22996 21732 23000 21788
rect 23000 21732 23056 21788
rect 23056 21732 23060 21788
rect 22996 21728 23060 21732
rect 23076 21788 23140 21792
rect 23076 21732 23080 21788
rect 23080 21732 23136 21788
rect 23136 21732 23140 21788
rect 23076 21728 23140 21732
rect 23156 21788 23220 21792
rect 23156 21732 23160 21788
rect 23160 21732 23216 21788
rect 23216 21732 23220 21788
rect 23156 21728 23220 21732
rect 23236 21788 23300 21792
rect 23236 21732 23240 21788
rect 23240 21732 23296 21788
rect 23296 21732 23300 21788
rect 23236 21728 23300 21732
rect 28916 21788 28980 21792
rect 28916 21732 28920 21788
rect 28920 21732 28976 21788
rect 28976 21732 28980 21788
rect 28916 21728 28980 21732
rect 28996 21788 29060 21792
rect 28996 21732 29000 21788
rect 29000 21732 29056 21788
rect 29056 21732 29060 21788
rect 28996 21728 29060 21732
rect 29076 21788 29140 21792
rect 29076 21732 29080 21788
rect 29080 21732 29136 21788
rect 29136 21732 29140 21788
rect 29076 21728 29140 21732
rect 29156 21788 29220 21792
rect 29156 21732 29160 21788
rect 29160 21732 29216 21788
rect 29216 21732 29220 21788
rect 29156 21728 29220 21732
rect 29236 21788 29300 21792
rect 29236 21732 29240 21788
rect 29240 21732 29296 21788
rect 29296 21732 29300 21788
rect 29236 21728 29300 21732
rect 4176 21244 4240 21248
rect 4176 21188 4180 21244
rect 4180 21188 4236 21244
rect 4236 21188 4240 21244
rect 4176 21184 4240 21188
rect 4256 21244 4320 21248
rect 4256 21188 4260 21244
rect 4260 21188 4316 21244
rect 4316 21188 4320 21244
rect 4256 21184 4320 21188
rect 4336 21244 4400 21248
rect 4336 21188 4340 21244
rect 4340 21188 4396 21244
rect 4396 21188 4400 21244
rect 4336 21184 4400 21188
rect 4416 21244 4480 21248
rect 4416 21188 4420 21244
rect 4420 21188 4476 21244
rect 4476 21188 4480 21244
rect 4416 21184 4480 21188
rect 4496 21244 4560 21248
rect 4496 21188 4500 21244
rect 4500 21188 4556 21244
rect 4556 21188 4560 21244
rect 4496 21184 4560 21188
rect 10176 21244 10240 21248
rect 10176 21188 10180 21244
rect 10180 21188 10236 21244
rect 10236 21188 10240 21244
rect 10176 21184 10240 21188
rect 10256 21244 10320 21248
rect 10256 21188 10260 21244
rect 10260 21188 10316 21244
rect 10316 21188 10320 21244
rect 10256 21184 10320 21188
rect 10336 21244 10400 21248
rect 10336 21188 10340 21244
rect 10340 21188 10396 21244
rect 10396 21188 10400 21244
rect 10336 21184 10400 21188
rect 10416 21244 10480 21248
rect 10416 21188 10420 21244
rect 10420 21188 10476 21244
rect 10476 21188 10480 21244
rect 10416 21184 10480 21188
rect 10496 21244 10560 21248
rect 10496 21188 10500 21244
rect 10500 21188 10556 21244
rect 10556 21188 10560 21244
rect 10496 21184 10560 21188
rect 16176 21244 16240 21248
rect 16176 21188 16180 21244
rect 16180 21188 16236 21244
rect 16236 21188 16240 21244
rect 16176 21184 16240 21188
rect 16256 21244 16320 21248
rect 16256 21188 16260 21244
rect 16260 21188 16316 21244
rect 16316 21188 16320 21244
rect 16256 21184 16320 21188
rect 16336 21244 16400 21248
rect 16336 21188 16340 21244
rect 16340 21188 16396 21244
rect 16396 21188 16400 21244
rect 16336 21184 16400 21188
rect 16416 21244 16480 21248
rect 16416 21188 16420 21244
rect 16420 21188 16476 21244
rect 16476 21188 16480 21244
rect 16416 21184 16480 21188
rect 16496 21244 16560 21248
rect 16496 21188 16500 21244
rect 16500 21188 16556 21244
rect 16556 21188 16560 21244
rect 16496 21184 16560 21188
rect 22176 21244 22240 21248
rect 22176 21188 22180 21244
rect 22180 21188 22236 21244
rect 22236 21188 22240 21244
rect 22176 21184 22240 21188
rect 22256 21244 22320 21248
rect 22256 21188 22260 21244
rect 22260 21188 22316 21244
rect 22316 21188 22320 21244
rect 22256 21184 22320 21188
rect 22336 21244 22400 21248
rect 22336 21188 22340 21244
rect 22340 21188 22396 21244
rect 22396 21188 22400 21244
rect 22336 21184 22400 21188
rect 22416 21244 22480 21248
rect 22416 21188 22420 21244
rect 22420 21188 22476 21244
rect 22476 21188 22480 21244
rect 22416 21184 22480 21188
rect 22496 21244 22560 21248
rect 22496 21188 22500 21244
rect 22500 21188 22556 21244
rect 22556 21188 22560 21244
rect 22496 21184 22560 21188
rect 28176 21244 28240 21248
rect 28176 21188 28180 21244
rect 28180 21188 28236 21244
rect 28236 21188 28240 21244
rect 28176 21184 28240 21188
rect 28256 21244 28320 21248
rect 28256 21188 28260 21244
rect 28260 21188 28316 21244
rect 28316 21188 28320 21244
rect 28256 21184 28320 21188
rect 28336 21244 28400 21248
rect 28336 21188 28340 21244
rect 28340 21188 28396 21244
rect 28396 21188 28400 21244
rect 28336 21184 28400 21188
rect 28416 21244 28480 21248
rect 28416 21188 28420 21244
rect 28420 21188 28476 21244
rect 28476 21188 28480 21244
rect 28416 21184 28480 21188
rect 28496 21244 28560 21248
rect 28496 21188 28500 21244
rect 28500 21188 28556 21244
rect 28556 21188 28560 21244
rect 28496 21184 28560 21188
rect 4916 20700 4980 20704
rect 4916 20644 4920 20700
rect 4920 20644 4976 20700
rect 4976 20644 4980 20700
rect 4916 20640 4980 20644
rect 4996 20700 5060 20704
rect 4996 20644 5000 20700
rect 5000 20644 5056 20700
rect 5056 20644 5060 20700
rect 4996 20640 5060 20644
rect 5076 20700 5140 20704
rect 5076 20644 5080 20700
rect 5080 20644 5136 20700
rect 5136 20644 5140 20700
rect 5076 20640 5140 20644
rect 5156 20700 5220 20704
rect 5156 20644 5160 20700
rect 5160 20644 5216 20700
rect 5216 20644 5220 20700
rect 5156 20640 5220 20644
rect 5236 20700 5300 20704
rect 5236 20644 5240 20700
rect 5240 20644 5296 20700
rect 5296 20644 5300 20700
rect 5236 20640 5300 20644
rect 10916 20700 10980 20704
rect 10916 20644 10920 20700
rect 10920 20644 10976 20700
rect 10976 20644 10980 20700
rect 10916 20640 10980 20644
rect 10996 20700 11060 20704
rect 10996 20644 11000 20700
rect 11000 20644 11056 20700
rect 11056 20644 11060 20700
rect 10996 20640 11060 20644
rect 11076 20700 11140 20704
rect 11076 20644 11080 20700
rect 11080 20644 11136 20700
rect 11136 20644 11140 20700
rect 11076 20640 11140 20644
rect 11156 20700 11220 20704
rect 11156 20644 11160 20700
rect 11160 20644 11216 20700
rect 11216 20644 11220 20700
rect 11156 20640 11220 20644
rect 11236 20700 11300 20704
rect 11236 20644 11240 20700
rect 11240 20644 11296 20700
rect 11296 20644 11300 20700
rect 11236 20640 11300 20644
rect 16916 20700 16980 20704
rect 16916 20644 16920 20700
rect 16920 20644 16976 20700
rect 16976 20644 16980 20700
rect 16916 20640 16980 20644
rect 16996 20700 17060 20704
rect 16996 20644 17000 20700
rect 17000 20644 17056 20700
rect 17056 20644 17060 20700
rect 16996 20640 17060 20644
rect 17076 20700 17140 20704
rect 17076 20644 17080 20700
rect 17080 20644 17136 20700
rect 17136 20644 17140 20700
rect 17076 20640 17140 20644
rect 17156 20700 17220 20704
rect 17156 20644 17160 20700
rect 17160 20644 17216 20700
rect 17216 20644 17220 20700
rect 17156 20640 17220 20644
rect 17236 20700 17300 20704
rect 17236 20644 17240 20700
rect 17240 20644 17296 20700
rect 17296 20644 17300 20700
rect 17236 20640 17300 20644
rect 22916 20700 22980 20704
rect 22916 20644 22920 20700
rect 22920 20644 22976 20700
rect 22976 20644 22980 20700
rect 22916 20640 22980 20644
rect 22996 20700 23060 20704
rect 22996 20644 23000 20700
rect 23000 20644 23056 20700
rect 23056 20644 23060 20700
rect 22996 20640 23060 20644
rect 23076 20700 23140 20704
rect 23076 20644 23080 20700
rect 23080 20644 23136 20700
rect 23136 20644 23140 20700
rect 23076 20640 23140 20644
rect 23156 20700 23220 20704
rect 23156 20644 23160 20700
rect 23160 20644 23216 20700
rect 23216 20644 23220 20700
rect 23156 20640 23220 20644
rect 23236 20700 23300 20704
rect 23236 20644 23240 20700
rect 23240 20644 23296 20700
rect 23296 20644 23300 20700
rect 23236 20640 23300 20644
rect 28916 20700 28980 20704
rect 28916 20644 28920 20700
rect 28920 20644 28976 20700
rect 28976 20644 28980 20700
rect 28916 20640 28980 20644
rect 28996 20700 29060 20704
rect 28996 20644 29000 20700
rect 29000 20644 29056 20700
rect 29056 20644 29060 20700
rect 28996 20640 29060 20644
rect 29076 20700 29140 20704
rect 29076 20644 29080 20700
rect 29080 20644 29136 20700
rect 29136 20644 29140 20700
rect 29076 20640 29140 20644
rect 29156 20700 29220 20704
rect 29156 20644 29160 20700
rect 29160 20644 29216 20700
rect 29216 20644 29220 20700
rect 29156 20640 29220 20644
rect 29236 20700 29300 20704
rect 29236 20644 29240 20700
rect 29240 20644 29296 20700
rect 29296 20644 29300 20700
rect 29236 20640 29300 20644
rect 4176 20156 4240 20160
rect 4176 20100 4180 20156
rect 4180 20100 4236 20156
rect 4236 20100 4240 20156
rect 4176 20096 4240 20100
rect 4256 20156 4320 20160
rect 4256 20100 4260 20156
rect 4260 20100 4316 20156
rect 4316 20100 4320 20156
rect 4256 20096 4320 20100
rect 4336 20156 4400 20160
rect 4336 20100 4340 20156
rect 4340 20100 4396 20156
rect 4396 20100 4400 20156
rect 4336 20096 4400 20100
rect 4416 20156 4480 20160
rect 4416 20100 4420 20156
rect 4420 20100 4476 20156
rect 4476 20100 4480 20156
rect 4416 20096 4480 20100
rect 4496 20156 4560 20160
rect 4496 20100 4500 20156
rect 4500 20100 4556 20156
rect 4556 20100 4560 20156
rect 4496 20096 4560 20100
rect 10176 20156 10240 20160
rect 10176 20100 10180 20156
rect 10180 20100 10236 20156
rect 10236 20100 10240 20156
rect 10176 20096 10240 20100
rect 10256 20156 10320 20160
rect 10256 20100 10260 20156
rect 10260 20100 10316 20156
rect 10316 20100 10320 20156
rect 10256 20096 10320 20100
rect 10336 20156 10400 20160
rect 10336 20100 10340 20156
rect 10340 20100 10396 20156
rect 10396 20100 10400 20156
rect 10336 20096 10400 20100
rect 10416 20156 10480 20160
rect 10416 20100 10420 20156
rect 10420 20100 10476 20156
rect 10476 20100 10480 20156
rect 10416 20096 10480 20100
rect 10496 20156 10560 20160
rect 10496 20100 10500 20156
rect 10500 20100 10556 20156
rect 10556 20100 10560 20156
rect 10496 20096 10560 20100
rect 16176 20156 16240 20160
rect 16176 20100 16180 20156
rect 16180 20100 16236 20156
rect 16236 20100 16240 20156
rect 16176 20096 16240 20100
rect 16256 20156 16320 20160
rect 16256 20100 16260 20156
rect 16260 20100 16316 20156
rect 16316 20100 16320 20156
rect 16256 20096 16320 20100
rect 16336 20156 16400 20160
rect 16336 20100 16340 20156
rect 16340 20100 16396 20156
rect 16396 20100 16400 20156
rect 16336 20096 16400 20100
rect 16416 20156 16480 20160
rect 16416 20100 16420 20156
rect 16420 20100 16476 20156
rect 16476 20100 16480 20156
rect 16416 20096 16480 20100
rect 16496 20156 16560 20160
rect 16496 20100 16500 20156
rect 16500 20100 16556 20156
rect 16556 20100 16560 20156
rect 16496 20096 16560 20100
rect 22176 20156 22240 20160
rect 22176 20100 22180 20156
rect 22180 20100 22236 20156
rect 22236 20100 22240 20156
rect 22176 20096 22240 20100
rect 22256 20156 22320 20160
rect 22256 20100 22260 20156
rect 22260 20100 22316 20156
rect 22316 20100 22320 20156
rect 22256 20096 22320 20100
rect 22336 20156 22400 20160
rect 22336 20100 22340 20156
rect 22340 20100 22396 20156
rect 22396 20100 22400 20156
rect 22336 20096 22400 20100
rect 22416 20156 22480 20160
rect 22416 20100 22420 20156
rect 22420 20100 22476 20156
rect 22476 20100 22480 20156
rect 22416 20096 22480 20100
rect 22496 20156 22560 20160
rect 22496 20100 22500 20156
rect 22500 20100 22556 20156
rect 22556 20100 22560 20156
rect 22496 20096 22560 20100
rect 28176 20156 28240 20160
rect 28176 20100 28180 20156
rect 28180 20100 28236 20156
rect 28236 20100 28240 20156
rect 28176 20096 28240 20100
rect 28256 20156 28320 20160
rect 28256 20100 28260 20156
rect 28260 20100 28316 20156
rect 28316 20100 28320 20156
rect 28256 20096 28320 20100
rect 28336 20156 28400 20160
rect 28336 20100 28340 20156
rect 28340 20100 28396 20156
rect 28396 20100 28400 20156
rect 28336 20096 28400 20100
rect 28416 20156 28480 20160
rect 28416 20100 28420 20156
rect 28420 20100 28476 20156
rect 28476 20100 28480 20156
rect 28416 20096 28480 20100
rect 28496 20156 28560 20160
rect 28496 20100 28500 20156
rect 28500 20100 28556 20156
rect 28556 20100 28560 20156
rect 28496 20096 28560 20100
rect 4916 19612 4980 19616
rect 4916 19556 4920 19612
rect 4920 19556 4976 19612
rect 4976 19556 4980 19612
rect 4916 19552 4980 19556
rect 4996 19612 5060 19616
rect 4996 19556 5000 19612
rect 5000 19556 5056 19612
rect 5056 19556 5060 19612
rect 4996 19552 5060 19556
rect 5076 19612 5140 19616
rect 5076 19556 5080 19612
rect 5080 19556 5136 19612
rect 5136 19556 5140 19612
rect 5076 19552 5140 19556
rect 5156 19612 5220 19616
rect 5156 19556 5160 19612
rect 5160 19556 5216 19612
rect 5216 19556 5220 19612
rect 5156 19552 5220 19556
rect 5236 19612 5300 19616
rect 5236 19556 5240 19612
rect 5240 19556 5296 19612
rect 5296 19556 5300 19612
rect 5236 19552 5300 19556
rect 10916 19612 10980 19616
rect 10916 19556 10920 19612
rect 10920 19556 10976 19612
rect 10976 19556 10980 19612
rect 10916 19552 10980 19556
rect 10996 19612 11060 19616
rect 10996 19556 11000 19612
rect 11000 19556 11056 19612
rect 11056 19556 11060 19612
rect 10996 19552 11060 19556
rect 11076 19612 11140 19616
rect 11076 19556 11080 19612
rect 11080 19556 11136 19612
rect 11136 19556 11140 19612
rect 11076 19552 11140 19556
rect 11156 19612 11220 19616
rect 11156 19556 11160 19612
rect 11160 19556 11216 19612
rect 11216 19556 11220 19612
rect 11156 19552 11220 19556
rect 11236 19612 11300 19616
rect 11236 19556 11240 19612
rect 11240 19556 11296 19612
rect 11296 19556 11300 19612
rect 11236 19552 11300 19556
rect 16916 19612 16980 19616
rect 16916 19556 16920 19612
rect 16920 19556 16976 19612
rect 16976 19556 16980 19612
rect 16916 19552 16980 19556
rect 16996 19612 17060 19616
rect 16996 19556 17000 19612
rect 17000 19556 17056 19612
rect 17056 19556 17060 19612
rect 16996 19552 17060 19556
rect 17076 19612 17140 19616
rect 17076 19556 17080 19612
rect 17080 19556 17136 19612
rect 17136 19556 17140 19612
rect 17076 19552 17140 19556
rect 17156 19612 17220 19616
rect 17156 19556 17160 19612
rect 17160 19556 17216 19612
rect 17216 19556 17220 19612
rect 17156 19552 17220 19556
rect 17236 19612 17300 19616
rect 17236 19556 17240 19612
rect 17240 19556 17296 19612
rect 17296 19556 17300 19612
rect 17236 19552 17300 19556
rect 22916 19612 22980 19616
rect 22916 19556 22920 19612
rect 22920 19556 22976 19612
rect 22976 19556 22980 19612
rect 22916 19552 22980 19556
rect 22996 19612 23060 19616
rect 22996 19556 23000 19612
rect 23000 19556 23056 19612
rect 23056 19556 23060 19612
rect 22996 19552 23060 19556
rect 23076 19612 23140 19616
rect 23076 19556 23080 19612
rect 23080 19556 23136 19612
rect 23136 19556 23140 19612
rect 23076 19552 23140 19556
rect 23156 19612 23220 19616
rect 23156 19556 23160 19612
rect 23160 19556 23216 19612
rect 23216 19556 23220 19612
rect 23156 19552 23220 19556
rect 23236 19612 23300 19616
rect 23236 19556 23240 19612
rect 23240 19556 23296 19612
rect 23296 19556 23300 19612
rect 23236 19552 23300 19556
rect 28916 19612 28980 19616
rect 28916 19556 28920 19612
rect 28920 19556 28976 19612
rect 28976 19556 28980 19612
rect 28916 19552 28980 19556
rect 28996 19612 29060 19616
rect 28996 19556 29000 19612
rect 29000 19556 29056 19612
rect 29056 19556 29060 19612
rect 28996 19552 29060 19556
rect 29076 19612 29140 19616
rect 29076 19556 29080 19612
rect 29080 19556 29136 19612
rect 29136 19556 29140 19612
rect 29076 19552 29140 19556
rect 29156 19612 29220 19616
rect 29156 19556 29160 19612
rect 29160 19556 29216 19612
rect 29216 19556 29220 19612
rect 29156 19552 29220 19556
rect 29236 19612 29300 19616
rect 29236 19556 29240 19612
rect 29240 19556 29296 19612
rect 29296 19556 29300 19612
rect 29236 19552 29300 19556
rect 4176 19068 4240 19072
rect 4176 19012 4180 19068
rect 4180 19012 4236 19068
rect 4236 19012 4240 19068
rect 4176 19008 4240 19012
rect 4256 19068 4320 19072
rect 4256 19012 4260 19068
rect 4260 19012 4316 19068
rect 4316 19012 4320 19068
rect 4256 19008 4320 19012
rect 4336 19068 4400 19072
rect 4336 19012 4340 19068
rect 4340 19012 4396 19068
rect 4396 19012 4400 19068
rect 4336 19008 4400 19012
rect 4416 19068 4480 19072
rect 4416 19012 4420 19068
rect 4420 19012 4476 19068
rect 4476 19012 4480 19068
rect 4416 19008 4480 19012
rect 4496 19068 4560 19072
rect 4496 19012 4500 19068
rect 4500 19012 4556 19068
rect 4556 19012 4560 19068
rect 4496 19008 4560 19012
rect 10176 19068 10240 19072
rect 10176 19012 10180 19068
rect 10180 19012 10236 19068
rect 10236 19012 10240 19068
rect 10176 19008 10240 19012
rect 10256 19068 10320 19072
rect 10256 19012 10260 19068
rect 10260 19012 10316 19068
rect 10316 19012 10320 19068
rect 10256 19008 10320 19012
rect 10336 19068 10400 19072
rect 10336 19012 10340 19068
rect 10340 19012 10396 19068
rect 10396 19012 10400 19068
rect 10336 19008 10400 19012
rect 10416 19068 10480 19072
rect 10416 19012 10420 19068
rect 10420 19012 10476 19068
rect 10476 19012 10480 19068
rect 10416 19008 10480 19012
rect 10496 19068 10560 19072
rect 10496 19012 10500 19068
rect 10500 19012 10556 19068
rect 10556 19012 10560 19068
rect 10496 19008 10560 19012
rect 16176 19068 16240 19072
rect 16176 19012 16180 19068
rect 16180 19012 16236 19068
rect 16236 19012 16240 19068
rect 16176 19008 16240 19012
rect 16256 19068 16320 19072
rect 16256 19012 16260 19068
rect 16260 19012 16316 19068
rect 16316 19012 16320 19068
rect 16256 19008 16320 19012
rect 16336 19068 16400 19072
rect 16336 19012 16340 19068
rect 16340 19012 16396 19068
rect 16396 19012 16400 19068
rect 16336 19008 16400 19012
rect 16416 19068 16480 19072
rect 16416 19012 16420 19068
rect 16420 19012 16476 19068
rect 16476 19012 16480 19068
rect 16416 19008 16480 19012
rect 16496 19068 16560 19072
rect 16496 19012 16500 19068
rect 16500 19012 16556 19068
rect 16556 19012 16560 19068
rect 16496 19008 16560 19012
rect 22176 19068 22240 19072
rect 22176 19012 22180 19068
rect 22180 19012 22236 19068
rect 22236 19012 22240 19068
rect 22176 19008 22240 19012
rect 22256 19068 22320 19072
rect 22256 19012 22260 19068
rect 22260 19012 22316 19068
rect 22316 19012 22320 19068
rect 22256 19008 22320 19012
rect 22336 19068 22400 19072
rect 22336 19012 22340 19068
rect 22340 19012 22396 19068
rect 22396 19012 22400 19068
rect 22336 19008 22400 19012
rect 22416 19068 22480 19072
rect 22416 19012 22420 19068
rect 22420 19012 22476 19068
rect 22476 19012 22480 19068
rect 22416 19008 22480 19012
rect 22496 19068 22560 19072
rect 22496 19012 22500 19068
rect 22500 19012 22556 19068
rect 22556 19012 22560 19068
rect 22496 19008 22560 19012
rect 28176 19068 28240 19072
rect 28176 19012 28180 19068
rect 28180 19012 28236 19068
rect 28236 19012 28240 19068
rect 28176 19008 28240 19012
rect 28256 19068 28320 19072
rect 28256 19012 28260 19068
rect 28260 19012 28316 19068
rect 28316 19012 28320 19068
rect 28256 19008 28320 19012
rect 28336 19068 28400 19072
rect 28336 19012 28340 19068
rect 28340 19012 28396 19068
rect 28396 19012 28400 19068
rect 28336 19008 28400 19012
rect 28416 19068 28480 19072
rect 28416 19012 28420 19068
rect 28420 19012 28476 19068
rect 28476 19012 28480 19068
rect 28416 19008 28480 19012
rect 28496 19068 28560 19072
rect 28496 19012 28500 19068
rect 28500 19012 28556 19068
rect 28556 19012 28560 19068
rect 28496 19008 28560 19012
rect 4916 18524 4980 18528
rect 4916 18468 4920 18524
rect 4920 18468 4976 18524
rect 4976 18468 4980 18524
rect 4916 18464 4980 18468
rect 4996 18524 5060 18528
rect 4996 18468 5000 18524
rect 5000 18468 5056 18524
rect 5056 18468 5060 18524
rect 4996 18464 5060 18468
rect 5076 18524 5140 18528
rect 5076 18468 5080 18524
rect 5080 18468 5136 18524
rect 5136 18468 5140 18524
rect 5076 18464 5140 18468
rect 5156 18524 5220 18528
rect 5156 18468 5160 18524
rect 5160 18468 5216 18524
rect 5216 18468 5220 18524
rect 5156 18464 5220 18468
rect 5236 18524 5300 18528
rect 5236 18468 5240 18524
rect 5240 18468 5296 18524
rect 5296 18468 5300 18524
rect 5236 18464 5300 18468
rect 10916 18524 10980 18528
rect 10916 18468 10920 18524
rect 10920 18468 10976 18524
rect 10976 18468 10980 18524
rect 10916 18464 10980 18468
rect 10996 18524 11060 18528
rect 10996 18468 11000 18524
rect 11000 18468 11056 18524
rect 11056 18468 11060 18524
rect 10996 18464 11060 18468
rect 11076 18524 11140 18528
rect 11076 18468 11080 18524
rect 11080 18468 11136 18524
rect 11136 18468 11140 18524
rect 11076 18464 11140 18468
rect 11156 18524 11220 18528
rect 11156 18468 11160 18524
rect 11160 18468 11216 18524
rect 11216 18468 11220 18524
rect 11156 18464 11220 18468
rect 11236 18524 11300 18528
rect 11236 18468 11240 18524
rect 11240 18468 11296 18524
rect 11296 18468 11300 18524
rect 11236 18464 11300 18468
rect 16916 18524 16980 18528
rect 16916 18468 16920 18524
rect 16920 18468 16976 18524
rect 16976 18468 16980 18524
rect 16916 18464 16980 18468
rect 16996 18524 17060 18528
rect 16996 18468 17000 18524
rect 17000 18468 17056 18524
rect 17056 18468 17060 18524
rect 16996 18464 17060 18468
rect 17076 18524 17140 18528
rect 17076 18468 17080 18524
rect 17080 18468 17136 18524
rect 17136 18468 17140 18524
rect 17076 18464 17140 18468
rect 17156 18524 17220 18528
rect 17156 18468 17160 18524
rect 17160 18468 17216 18524
rect 17216 18468 17220 18524
rect 17156 18464 17220 18468
rect 17236 18524 17300 18528
rect 17236 18468 17240 18524
rect 17240 18468 17296 18524
rect 17296 18468 17300 18524
rect 17236 18464 17300 18468
rect 22916 18524 22980 18528
rect 22916 18468 22920 18524
rect 22920 18468 22976 18524
rect 22976 18468 22980 18524
rect 22916 18464 22980 18468
rect 22996 18524 23060 18528
rect 22996 18468 23000 18524
rect 23000 18468 23056 18524
rect 23056 18468 23060 18524
rect 22996 18464 23060 18468
rect 23076 18524 23140 18528
rect 23076 18468 23080 18524
rect 23080 18468 23136 18524
rect 23136 18468 23140 18524
rect 23076 18464 23140 18468
rect 23156 18524 23220 18528
rect 23156 18468 23160 18524
rect 23160 18468 23216 18524
rect 23216 18468 23220 18524
rect 23156 18464 23220 18468
rect 23236 18524 23300 18528
rect 23236 18468 23240 18524
rect 23240 18468 23296 18524
rect 23296 18468 23300 18524
rect 23236 18464 23300 18468
rect 28916 18524 28980 18528
rect 28916 18468 28920 18524
rect 28920 18468 28976 18524
rect 28976 18468 28980 18524
rect 28916 18464 28980 18468
rect 28996 18524 29060 18528
rect 28996 18468 29000 18524
rect 29000 18468 29056 18524
rect 29056 18468 29060 18524
rect 28996 18464 29060 18468
rect 29076 18524 29140 18528
rect 29076 18468 29080 18524
rect 29080 18468 29136 18524
rect 29136 18468 29140 18524
rect 29076 18464 29140 18468
rect 29156 18524 29220 18528
rect 29156 18468 29160 18524
rect 29160 18468 29216 18524
rect 29216 18468 29220 18524
rect 29156 18464 29220 18468
rect 29236 18524 29300 18528
rect 29236 18468 29240 18524
rect 29240 18468 29296 18524
rect 29296 18468 29300 18524
rect 29236 18464 29300 18468
rect 4176 17980 4240 17984
rect 4176 17924 4180 17980
rect 4180 17924 4236 17980
rect 4236 17924 4240 17980
rect 4176 17920 4240 17924
rect 4256 17980 4320 17984
rect 4256 17924 4260 17980
rect 4260 17924 4316 17980
rect 4316 17924 4320 17980
rect 4256 17920 4320 17924
rect 4336 17980 4400 17984
rect 4336 17924 4340 17980
rect 4340 17924 4396 17980
rect 4396 17924 4400 17980
rect 4336 17920 4400 17924
rect 4416 17980 4480 17984
rect 4416 17924 4420 17980
rect 4420 17924 4476 17980
rect 4476 17924 4480 17980
rect 4416 17920 4480 17924
rect 4496 17980 4560 17984
rect 4496 17924 4500 17980
rect 4500 17924 4556 17980
rect 4556 17924 4560 17980
rect 4496 17920 4560 17924
rect 10176 17980 10240 17984
rect 10176 17924 10180 17980
rect 10180 17924 10236 17980
rect 10236 17924 10240 17980
rect 10176 17920 10240 17924
rect 10256 17980 10320 17984
rect 10256 17924 10260 17980
rect 10260 17924 10316 17980
rect 10316 17924 10320 17980
rect 10256 17920 10320 17924
rect 10336 17980 10400 17984
rect 10336 17924 10340 17980
rect 10340 17924 10396 17980
rect 10396 17924 10400 17980
rect 10336 17920 10400 17924
rect 10416 17980 10480 17984
rect 10416 17924 10420 17980
rect 10420 17924 10476 17980
rect 10476 17924 10480 17980
rect 10416 17920 10480 17924
rect 10496 17980 10560 17984
rect 10496 17924 10500 17980
rect 10500 17924 10556 17980
rect 10556 17924 10560 17980
rect 10496 17920 10560 17924
rect 16176 17980 16240 17984
rect 16176 17924 16180 17980
rect 16180 17924 16236 17980
rect 16236 17924 16240 17980
rect 16176 17920 16240 17924
rect 16256 17980 16320 17984
rect 16256 17924 16260 17980
rect 16260 17924 16316 17980
rect 16316 17924 16320 17980
rect 16256 17920 16320 17924
rect 16336 17980 16400 17984
rect 16336 17924 16340 17980
rect 16340 17924 16396 17980
rect 16396 17924 16400 17980
rect 16336 17920 16400 17924
rect 16416 17980 16480 17984
rect 16416 17924 16420 17980
rect 16420 17924 16476 17980
rect 16476 17924 16480 17980
rect 16416 17920 16480 17924
rect 16496 17980 16560 17984
rect 16496 17924 16500 17980
rect 16500 17924 16556 17980
rect 16556 17924 16560 17980
rect 16496 17920 16560 17924
rect 22176 17980 22240 17984
rect 22176 17924 22180 17980
rect 22180 17924 22236 17980
rect 22236 17924 22240 17980
rect 22176 17920 22240 17924
rect 22256 17980 22320 17984
rect 22256 17924 22260 17980
rect 22260 17924 22316 17980
rect 22316 17924 22320 17980
rect 22256 17920 22320 17924
rect 22336 17980 22400 17984
rect 22336 17924 22340 17980
rect 22340 17924 22396 17980
rect 22396 17924 22400 17980
rect 22336 17920 22400 17924
rect 22416 17980 22480 17984
rect 22416 17924 22420 17980
rect 22420 17924 22476 17980
rect 22476 17924 22480 17980
rect 22416 17920 22480 17924
rect 22496 17980 22560 17984
rect 22496 17924 22500 17980
rect 22500 17924 22556 17980
rect 22556 17924 22560 17980
rect 22496 17920 22560 17924
rect 28176 17980 28240 17984
rect 28176 17924 28180 17980
rect 28180 17924 28236 17980
rect 28236 17924 28240 17980
rect 28176 17920 28240 17924
rect 28256 17980 28320 17984
rect 28256 17924 28260 17980
rect 28260 17924 28316 17980
rect 28316 17924 28320 17980
rect 28256 17920 28320 17924
rect 28336 17980 28400 17984
rect 28336 17924 28340 17980
rect 28340 17924 28396 17980
rect 28396 17924 28400 17980
rect 28336 17920 28400 17924
rect 28416 17980 28480 17984
rect 28416 17924 28420 17980
rect 28420 17924 28476 17980
rect 28476 17924 28480 17980
rect 28416 17920 28480 17924
rect 28496 17980 28560 17984
rect 28496 17924 28500 17980
rect 28500 17924 28556 17980
rect 28556 17924 28560 17980
rect 28496 17920 28560 17924
rect 4916 17436 4980 17440
rect 4916 17380 4920 17436
rect 4920 17380 4976 17436
rect 4976 17380 4980 17436
rect 4916 17376 4980 17380
rect 4996 17436 5060 17440
rect 4996 17380 5000 17436
rect 5000 17380 5056 17436
rect 5056 17380 5060 17436
rect 4996 17376 5060 17380
rect 5076 17436 5140 17440
rect 5076 17380 5080 17436
rect 5080 17380 5136 17436
rect 5136 17380 5140 17436
rect 5076 17376 5140 17380
rect 5156 17436 5220 17440
rect 5156 17380 5160 17436
rect 5160 17380 5216 17436
rect 5216 17380 5220 17436
rect 5156 17376 5220 17380
rect 5236 17436 5300 17440
rect 5236 17380 5240 17436
rect 5240 17380 5296 17436
rect 5296 17380 5300 17436
rect 5236 17376 5300 17380
rect 10916 17436 10980 17440
rect 10916 17380 10920 17436
rect 10920 17380 10976 17436
rect 10976 17380 10980 17436
rect 10916 17376 10980 17380
rect 10996 17436 11060 17440
rect 10996 17380 11000 17436
rect 11000 17380 11056 17436
rect 11056 17380 11060 17436
rect 10996 17376 11060 17380
rect 11076 17436 11140 17440
rect 11076 17380 11080 17436
rect 11080 17380 11136 17436
rect 11136 17380 11140 17436
rect 11076 17376 11140 17380
rect 11156 17436 11220 17440
rect 11156 17380 11160 17436
rect 11160 17380 11216 17436
rect 11216 17380 11220 17436
rect 11156 17376 11220 17380
rect 11236 17436 11300 17440
rect 11236 17380 11240 17436
rect 11240 17380 11296 17436
rect 11296 17380 11300 17436
rect 11236 17376 11300 17380
rect 16916 17436 16980 17440
rect 16916 17380 16920 17436
rect 16920 17380 16976 17436
rect 16976 17380 16980 17436
rect 16916 17376 16980 17380
rect 16996 17436 17060 17440
rect 16996 17380 17000 17436
rect 17000 17380 17056 17436
rect 17056 17380 17060 17436
rect 16996 17376 17060 17380
rect 17076 17436 17140 17440
rect 17076 17380 17080 17436
rect 17080 17380 17136 17436
rect 17136 17380 17140 17436
rect 17076 17376 17140 17380
rect 17156 17436 17220 17440
rect 17156 17380 17160 17436
rect 17160 17380 17216 17436
rect 17216 17380 17220 17436
rect 17156 17376 17220 17380
rect 17236 17436 17300 17440
rect 17236 17380 17240 17436
rect 17240 17380 17296 17436
rect 17296 17380 17300 17436
rect 17236 17376 17300 17380
rect 22916 17436 22980 17440
rect 22916 17380 22920 17436
rect 22920 17380 22976 17436
rect 22976 17380 22980 17436
rect 22916 17376 22980 17380
rect 22996 17436 23060 17440
rect 22996 17380 23000 17436
rect 23000 17380 23056 17436
rect 23056 17380 23060 17436
rect 22996 17376 23060 17380
rect 23076 17436 23140 17440
rect 23076 17380 23080 17436
rect 23080 17380 23136 17436
rect 23136 17380 23140 17436
rect 23076 17376 23140 17380
rect 23156 17436 23220 17440
rect 23156 17380 23160 17436
rect 23160 17380 23216 17436
rect 23216 17380 23220 17436
rect 23156 17376 23220 17380
rect 23236 17436 23300 17440
rect 23236 17380 23240 17436
rect 23240 17380 23296 17436
rect 23296 17380 23300 17436
rect 23236 17376 23300 17380
rect 28916 17436 28980 17440
rect 28916 17380 28920 17436
rect 28920 17380 28976 17436
rect 28976 17380 28980 17436
rect 28916 17376 28980 17380
rect 28996 17436 29060 17440
rect 28996 17380 29000 17436
rect 29000 17380 29056 17436
rect 29056 17380 29060 17436
rect 28996 17376 29060 17380
rect 29076 17436 29140 17440
rect 29076 17380 29080 17436
rect 29080 17380 29136 17436
rect 29136 17380 29140 17436
rect 29076 17376 29140 17380
rect 29156 17436 29220 17440
rect 29156 17380 29160 17436
rect 29160 17380 29216 17436
rect 29216 17380 29220 17436
rect 29156 17376 29220 17380
rect 29236 17436 29300 17440
rect 29236 17380 29240 17436
rect 29240 17380 29296 17436
rect 29296 17380 29300 17436
rect 29236 17376 29300 17380
rect 15332 17308 15396 17372
rect 27844 17172 27908 17236
rect 4176 16892 4240 16896
rect 4176 16836 4180 16892
rect 4180 16836 4236 16892
rect 4236 16836 4240 16892
rect 4176 16832 4240 16836
rect 4256 16892 4320 16896
rect 4256 16836 4260 16892
rect 4260 16836 4316 16892
rect 4316 16836 4320 16892
rect 4256 16832 4320 16836
rect 4336 16892 4400 16896
rect 4336 16836 4340 16892
rect 4340 16836 4396 16892
rect 4396 16836 4400 16892
rect 4336 16832 4400 16836
rect 4416 16892 4480 16896
rect 4416 16836 4420 16892
rect 4420 16836 4476 16892
rect 4476 16836 4480 16892
rect 4416 16832 4480 16836
rect 4496 16892 4560 16896
rect 4496 16836 4500 16892
rect 4500 16836 4556 16892
rect 4556 16836 4560 16892
rect 4496 16832 4560 16836
rect 10176 16892 10240 16896
rect 10176 16836 10180 16892
rect 10180 16836 10236 16892
rect 10236 16836 10240 16892
rect 10176 16832 10240 16836
rect 10256 16892 10320 16896
rect 10256 16836 10260 16892
rect 10260 16836 10316 16892
rect 10316 16836 10320 16892
rect 10256 16832 10320 16836
rect 10336 16892 10400 16896
rect 10336 16836 10340 16892
rect 10340 16836 10396 16892
rect 10396 16836 10400 16892
rect 10336 16832 10400 16836
rect 10416 16892 10480 16896
rect 10416 16836 10420 16892
rect 10420 16836 10476 16892
rect 10476 16836 10480 16892
rect 10416 16832 10480 16836
rect 10496 16892 10560 16896
rect 10496 16836 10500 16892
rect 10500 16836 10556 16892
rect 10556 16836 10560 16892
rect 10496 16832 10560 16836
rect 16176 16892 16240 16896
rect 16176 16836 16180 16892
rect 16180 16836 16236 16892
rect 16236 16836 16240 16892
rect 16176 16832 16240 16836
rect 16256 16892 16320 16896
rect 16256 16836 16260 16892
rect 16260 16836 16316 16892
rect 16316 16836 16320 16892
rect 16256 16832 16320 16836
rect 16336 16892 16400 16896
rect 16336 16836 16340 16892
rect 16340 16836 16396 16892
rect 16396 16836 16400 16892
rect 16336 16832 16400 16836
rect 16416 16892 16480 16896
rect 16416 16836 16420 16892
rect 16420 16836 16476 16892
rect 16476 16836 16480 16892
rect 16416 16832 16480 16836
rect 16496 16892 16560 16896
rect 16496 16836 16500 16892
rect 16500 16836 16556 16892
rect 16556 16836 16560 16892
rect 16496 16832 16560 16836
rect 22176 16892 22240 16896
rect 22176 16836 22180 16892
rect 22180 16836 22236 16892
rect 22236 16836 22240 16892
rect 22176 16832 22240 16836
rect 22256 16892 22320 16896
rect 22256 16836 22260 16892
rect 22260 16836 22316 16892
rect 22316 16836 22320 16892
rect 22256 16832 22320 16836
rect 22336 16892 22400 16896
rect 22336 16836 22340 16892
rect 22340 16836 22396 16892
rect 22396 16836 22400 16892
rect 22336 16832 22400 16836
rect 22416 16892 22480 16896
rect 22416 16836 22420 16892
rect 22420 16836 22476 16892
rect 22476 16836 22480 16892
rect 22416 16832 22480 16836
rect 22496 16892 22560 16896
rect 22496 16836 22500 16892
rect 22500 16836 22556 16892
rect 22556 16836 22560 16892
rect 22496 16832 22560 16836
rect 28176 16892 28240 16896
rect 28176 16836 28180 16892
rect 28180 16836 28236 16892
rect 28236 16836 28240 16892
rect 28176 16832 28240 16836
rect 28256 16892 28320 16896
rect 28256 16836 28260 16892
rect 28260 16836 28316 16892
rect 28316 16836 28320 16892
rect 28256 16832 28320 16836
rect 28336 16892 28400 16896
rect 28336 16836 28340 16892
rect 28340 16836 28396 16892
rect 28396 16836 28400 16892
rect 28336 16832 28400 16836
rect 28416 16892 28480 16896
rect 28416 16836 28420 16892
rect 28420 16836 28476 16892
rect 28476 16836 28480 16892
rect 28416 16832 28480 16836
rect 28496 16892 28560 16896
rect 28496 16836 28500 16892
rect 28500 16836 28556 16892
rect 28556 16836 28560 16892
rect 28496 16832 28560 16836
rect 4916 16348 4980 16352
rect 4916 16292 4920 16348
rect 4920 16292 4976 16348
rect 4976 16292 4980 16348
rect 4916 16288 4980 16292
rect 4996 16348 5060 16352
rect 4996 16292 5000 16348
rect 5000 16292 5056 16348
rect 5056 16292 5060 16348
rect 4996 16288 5060 16292
rect 5076 16348 5140 16352
rect 5076 16292 5080 16348
rect 5080 16292 5136 16348
rect 5136 16292 5140 16348
rect 5076 16288 5140 16292
rect 5156 16348 5220 16352
rect 5156 16292 5160 16348
rect 5160 16292 5216 16348
rect 5216 16292 5220 16348
rect 5156 16288 5220 16292
rect 5236 16348 5300 16352
rect 5236 16292 5240 16348
rect 5240 16292 5296 16348
rect 5296 16292 5300 16348
rect 5236 16288 5300 16292
rect 10916 16348 10980 16352
rect 10916 16292 10920 16348
rect 10920 16292 10976 16348
rect 10976 16292 10980 16348
rect 10916 16288 10980 16292
rect 10996 16348 11060 16352
rect 10996 16292 11000 16348
rect 11000 16292 11056 16348
rect 11056 16292 11060 16348
rect 10996 16288 11060 16292
rect 11076 16348 11140 16352
rect 11076 16292 11080 16348
rect 11080 16292 11136 16348
rect 11136 16292 11140 16348
rect 11076 16288 11140 16292
rect 11156 16348 11220 16352
rect 11156 16292 11160 16348
rect 11160 16292 11216 16348
rect 11216 16292 11220 16348
rect 11156 16288 11220 16292
rect 11236 16348 11300 16352
rect 11236 16292 11240 16348
rect 11240 16292 11296 16348
rect 11296 16292 11300 16348
rect 11236 16288 11300 16292
rect 16916 16348 16980 16352
rect 16916 16292 16920 16348
rect 16920 16292 16976 16348
rect 16976 16292 16980 16348
rect 16916 16288 16980 16292
rect 16996 16348 17060 16352
rect 16996 16292 17000 16348
rect 17000 16292 17056 16348
rect 17056 16292 17060 16348
rect 16996 16288 17060 16292
rect 17076 16348 17140 16352
rect 17076 16292 17080 16348
rect 17080 16292 17136 16348
rect 17136 16292 17140 16348
rect 17076 16288 17140 16292
rect 17156 16348 17220 16352
rect 17156 16292 17160 16348
rect 17160 16292 17216 16348
rect 17216 16292 17220 16348
rect 17156 16288 17220 16292
rect 17236 16348 17300 16352
rect 17236 16292 17240 16348
rect 17240 16292 17296 16348
rect 17296 16292 17300 16348
rect 17236 16288 17300 16292
rect 22916 16348 22980 16352
rect 22916 16292 22920 16348
rect 22920 16292 22976 16348
rect 22976 16292 22980 16348
rect 22916 16288 22980 16292
rect 22996 16348 23060 16352
rect 22996 16292 23000 16348
rect 23000 16292 23056 16348
rect 23056 16292 23060 16348
rect 22996 16288 23060 16292
rect 23076 16348 23140 16352
rect 23076 16292 23080 16348
rect 23080 16292 23136 16348
rect 23136 16292 23140 16348
rect 23076 16288 23140 16292
rect 23156 16348 23220 16352
rect 23156 16292 23160 16348
rect 23160 16292 23216 16348
rect 23216 16292 23220 16348
rect 23156 16288 23220 16292
rect 23236 16348 23300 16352
rect 23236 16292 23240 16348
rect 23240 16292 23296 16348
rect 23296 16292 23300 16348
rect 23236 16288 23300 16292
rect 28916 16348 28980 16352
rect 28916 16292 28920 16348
rect 28920 16292 28976 16348
rect 28976 16292 28980 16348
rect 28916 16288 28980 16292
rect 28996 16348 29060 16352
rect 28996 16292 29000 16348
rect 29000 16292 29056 16348
rect 29056 16292 29060 16348
rect 28996 16288 29060 16292
rect 29076 16348 29140 16352
rect 29076 16292 29080 16348
rect 29080 16292 29136 16348
rect 29136 16292 29140 16348
rect 29076 16288 29140 16292
rect 29156 16348 29220 16352
rect 29156 16292 29160 16348
rect 29160 16292 29216 16348
rect 29216 16292 29220 16348
rect 29156 16288 29220 16292
rect 29236 16348 29300 16352
rect 29236 16292 29240 16348
rect 29240 16292 29296 16348
rect 29296 16292 29300 16348
rect 29236 16288 29300 16292
rect 4176 15804 4240 15808
rect 4176 15748 4180 15804
rect 4180 15748 4236 15804
rect 4236 15748 4240 15804
rect 4176 15744 4240 15748
rect 4256 15804 4320 15808
rect 4256 15748 4260 15804
rect 4260 15748 4316 15804
rect 4316 15748 4320 15804
rect 4256 15744 4320 15748
rect 4336 15804 4400 15808
rect 4336 15748 4340 15804
rect 4340 15748 4396 15804
rect 4396 15748 4400 15804
rect 4336 15744 4400 15748
rect 4416 15804 4480 15808
rect 4416 15748 4420 15804
rect 4420 15748 4476 15804
rect 4476 15748 4480 15804
rect 4416 15744 4480 15748
rect 4496 15804 4560 15808
rect 4496 15748 4500 15804
rect 4500 15748 4556 15804
rect 4556 15748 4560 15804
rect 4496 15744 4560 15748
rect 10176 15804 10240 15808
rect 10176 15748 10180 15804
rect 10180 15748 10236 15804
rect 10236 15748 10240 15804
rect 10176 15744 10240 15748
rect 10256 15804 10320 15808
rect 10256 15748 10260 15804
rect 10260 15748 10316 15804
rect 10316 15748 10320 15804
rect 10256 15744 10320 15748
rect 10336 15804 10400 15808
rect 10336 15748 10340 15804
rect 10340 15748 10396 15804
rect 10396 15748 10400 15804
rect 10336 15744 10400 15748
rect 10416 15804 10480 15808
rect 10416 15748 10420 15804
rect 10420 15748 10476 15804
rect 10476 15748 10480 15804
rect 10416 15744 10480 15748
rect 10496 15804 10560 15808
rect 10496 15748 10500 15804
rect 10500 15748 10556 15804
rect 10556 15748 10560 15804
rect 10496 15744 10560 15748
rect 16176 15804 16240 15808
rect 16176 15748 16180 15804
rect 16180 15748 16236 15804
rect 16236 15748 16240 15804
rect 16176 15744 16240 15748
rect 16256 15804 16320 15808
rect 16256 15748 16260 15804
rect 16260 15748 16316 15804
rect 16316 15748 16320 15804
rect 16256 15744 16320 15748
rect 16336 15804 16400 15808
rect 16336 15748 16340 15804
rect 16340 15748 16396 15804
rect 16396 15748 16400 15804
rect 16336 15744 16400 15748
rect 16416 15804 16480 15808
rect 16416 15748 16420 15804
rect 16420 15748 16476 15804
rect 16476 15748 16480 15804
rect 16416 15744 16480 15748
rect 16496 15804 16560 15808
rect 16496 15748 16500 15804
rect 16500 15748 16556 15804
rect 16556 15748 16560 15804
rect 16496 15744 16560 15748
rect 22176 15804 22240 15808
rect 22176 15748 22180 15804
rect 22180 15748 22236 15804
rect 22236 15748 22240 15804
rect 22176 15744 22240 15748
rect 22256 15804 22320 15808
rect 22256 15748 22260 15804
rect 22260 15748 22316 15804
rect 22316 15748 22320 15804
rect 22256 15744 22320 15748
rect 22336 15804 22400 15808
rect 22336 15748 22340 15804
rect 22340 15748 22396 15804
rect 22396 15748 22400 15804
rect 22336 15744 22400 15748
rect 22416 15804 22480 15808
rect 22416 15748 22420 15804
rect 22420 15748 22476 15804
rect 22476 15748 22480 15804
rect 22416 15744 22480 15748
rect 22496 15804 22560 15808
rect 22496 15748 22500 15804
rect 22500 15748 22556 15804
rect 22556 15748 22560 15804
rect 22496 15744 22560 15748
rect 28176 15804 28240 15808
rect 28176 15748 28180 15804
rect 28180 15748 28236 15804
rect 28236 15748 28240 15804
rect 28176 15744 28240 15748
rect 28256 15804 28320 15808
rect 28256 15748 28260 15804
rect 28260 15748 28316 15804
rect 28316 15748 28320 15804
rect 28256 15744 28320 15748
rect 28336 15804 28400 15808
rect 28336 15748 28340 15804
rect 28340 15748 28396 15804
rect 28396 15748 28400 15804
rect 28336 15744 28400 15748
rect 28416 15804 28480 15808
rect 28416 15748 28420 15804
rect 28420 15748 28476 15804
rect 28476 15748 28480 15804
rect 28416 15744 28480 15748
rect 28496 15804 28560 15808
rect 28496 15748 28500 15804
rect 28500 15748 28556 15804
rect 28556 15748 28560 15804
rect 28496 15744 28560 15748
rect 4916 15260 4980 15264
rect 4916 15204 4920 15260
rect 4920 15204 4976 15260
rect 4976 15204 4980 15260
rect 4916 15200 4980 15204
rect 4996 15260 5060 15264
rect 4996 15204 5000 15260
rect 5000 15204 5056 15260
rect 5056 15204 5060 15260
rect 4996 15200 5060 15204
rect 5076 15260 5140 15264
rect 5076 15204 5080 15260
rect 5080 15204 5136 15260
rect 5136 15204 5140 15260
rect 5076 15200 5140 15204
rect 5156 15260 5220 15264
rect 5156 15204 5160 15260
rect 5160 15204 5216 15260
rect 5216 15204 5220 15260
rect 5156 15200 5220 15204
rect 5236 15260 5300 15264
rect 5236 15204 5240 15260
rect 5240 15204 5296 15260
rect 5296 15204 5300 15260
rect 5236 15200 5300 15204
rect 10916 15260 10980 15264
rect 10916 15204 10920 15260
rect 10920 15204 10976 15260
rect 10976 15204 10980 15260
rect 10916 15200 10980 15204
rect 10996 15260 11060 15264
rect 10996 15204 11000 15260
rect 11000 15204 11056 15260
rect 11056 15204 11060 15260
rect 10996 15200 11060 15204
rect 11076 15260 11140 15264
rect 11076 15204 11080 15260
rect 11080 15204 11136 15260
rect 11136 15204 11140 15260
rect 11076 15200 11140 15204
rect 11156 15260 11220 15264
rect 11156 15204 11160 15260
rect 11160 15204 11216 15260
rect 11216 15204 11220 15260
rect 11156 15200 11220 15204
rect 11236 15260 11300 15264
rect 11236 15204 11240 15260
rect 11240 15204 11296 15260
rect 11296 15204 11300 15260
rect 11236 15200 11300 15204
rect 16916 15260 16980 15264
rect 16916 15204 16920 15260
rect 16920 15204 16976 15260
rect 16976 15204 16980 15260
rect 16916 15200 16980 15204
rect 16996 15260 17060 15264
rect 16996 15204 17000 15260
rect 17000 15204 17056 15260
rect 17056 15204 17060 15260
rect 16996 15200 17060 15204
rect 17076 15260 17140 15264
rect 17076 15204 17080 15260
rect 17080 15204 17136 15260
rect 17136 15204 17140 15260
rect 17076 15200 17140 15204
rect 17156 15260 17220 15264
rect 17156 15204 17160 15260
rect 17160 15204 17216 15260
rect 17216 15204 17220 15260
rect 17156 15200 17220 15204
rect 17236 15260 17300 15264
rect 17236 15204 17240 15260
rect 17240 15204 17296 15260
rect 17296 15204 17300 15260
rect 17236 15200 17300 15204
rect 22916 15260 22980 15264
rect 22916 15204 22920 15260
rect 22920 15204 22976 15260
rect 22976 15204 22980 15260
rect 22916 15200 22980 15204
rect 22996 15260 23060 15264
rect 22996 15204 23000 15260
rect 23000 15204 23056 15260
rect 23056 15204 23060 15260
rect 22996 15200 23060 15204
rect 23076 15260 23140 15264
rect 23076 15204 23080 15260
rect 23080 15204 23136 15260
rect 23136 15204 23140 15260
rect 23076 15200 23140 15204
rect 23156 15260 23220 15264
rect 23156 15204 23160 15260
rect 23160 15204 23216 15260
rect 23216 15204 23220 15260
rect 23156 15200 23220 15204
rect 23236 15260 23300 15264
rect 23236 15204 23240 15260
rect 23240 15204 23296 15260
rect 23296 15204 23300 15260
rect 23236 15200 23300 15204
rect 28916 15260 28980 15264
rect 28916 15204 28920 15260
rect 28920 15204 28976 15260
rect 28976 15204 28980 15260
rect 28916 15200 28980 15204
rect 28996 15260 29060 15264
rect 28996 15204 29000 15260
rect 29000 15204 29056 15260
rect 29056 15204 29060 15260
rect 28996 15200 29060 15204
rect 29076 15260 29140 15264
rect 29076 15204 29080 15260
rect 29080 15204 29136 15260
rect 29136 15204 29140 15260
rect 29076 15200 29140 15204
rect 29156 15260 29220 15264
rect 29156 15204 29160 15260
rect 29160 15204 29216 15260
rect 29216 15204 29220 15260
rect 29156 15200 29220 15204
rect 29236 15260 29300 15264
rect 29236 15204 29240 15260
rect 29240 15204 29296 15260
rect 29296 15204 29300 15260
rect 29236 15200 29300 15204
rect 24532 15132 24596 15196
rect 4176 14716 4240 14720
rect 4176 14660 4180 14716
rect 4180 14660 4236 14716
rect 4236 14660 4240 14716
rect 4176 14656 4240 14660
rect 4256 14716 4320 14720
rect 4256 14660 4260 14716
rect 4260 14660 4316 14716
rect 4316 14660 4320 14716
rect 4256 14656 4320 14660
rect 4336 14716 4400 14720
rect 4336 14660 4340 14716
rect 4340 14660 4396 14716
rect 4396 14660 4400 14716
rect 4336 14656 4400 14660
rect 4416 14716 4480 14720
rect 4416 14660 4420 14716
rect 4420 14660 4476 14716
rect 4476 14660 4480 14716
rect 4416 14656 4480 14660
rect 4496 14716 4560 14720
rect 4496 14660 4500 14716
rect 4500 14660 4556 14716
rect 4556 14660 4560 14716
rect 4496 14656 4560 14660
rect 10176 14716 10240 14720
rect 10176 14660 10180 14716
rect 10180 14660 10236 14716
rect 10236 14660 10240 14716
rect 10176 14656 10240 14660
rect 10256 14716 10320 14720
rect 10256 14660 10260 14716
rect 10260 14660 10316 14716
rect 10316 14660 10320 14716
rect 10256 14656 10320 14660
rect 10336 14716 10400 14720
rect 10336 14660 10340 14716
rect 10340 14660 10396 14716
rect 10396 14660 10400 14716
rect 10336 14656 10400 14660
rect 10416 14716 10480 14720
rect 10416 14660 10420 14716
rect 10420 14660 10476 14716
rect 10476 14660 10480 14716
rect 10416 14656 10480 14660
rect 10496 14716 10560 14720
rect 10496 14660 10500 14716
rect 10500 14660 10556 14716
rect 10556 14660 10560 14716
rect 10496 14656 10560 14660
rect 16176 14716 16240 14720
rect 16176 14660 16180 14716
rect 16180 14660 16236 14716
rect 16236 14660 16240 14716
rect 16176 14656 16240 14660
rect 16256 14716 16320 14720
rect 16256 14660 16260 14716
rect 16260 14660 16316 14716
rect 16316 14660 16320 14716
rect 16256 14656 16320 14660
rect 16336 14716 16400 14720
rect 16336 14660 16340 14716
rect 16340 14660 16396 14716
rect 16396 14660 16400 14716
rect 16336 14656 16400 14660
rect 16416 14716 16480 14720
rect 16416 14660 16420 14716
rect 16420 14660 16476 14716
rect 16476 14660 16480 14716
rect 16416 14656 16480 14660
rect 16496 14716 16560 14720
rect 16496 14660 16500 14716
rect 16500 14660 16556 14716
rect 16556 14660 16560 14716
rect 16496 14656 16560 14660
rect 22176 14716 22240 14720
rect 22176 14660 22180 14716
rect 22180 14660 22236 14716
rect 22236 14660 22240 14716
rect 22176 14656 22240 14660
rect 22256 14716 22320 14720
rect 22256 14660 22260 14716
rect 22260 14660 22316 14716
rect 22316 14660 22320 14716
rect 22256 14656 22320 14660
rect 22336 14716 22400 14720
rect 22336 14660 22340 14716
rect 22340 14660 22396 14716
rect 22396 14660 22400 14716
rect 22336 14656 22400 14660
rect 22416 14716 22480 14720
rect 22416 14660 22420 14716
rect 22420 14660 22476 14716
rect 22476 14660 22480 14716
rect 22416 14656 22480 14660
rect 22496 14716 22560 14720
rect 22496 14660 22500 14716
rect 22500 14660 22556 14716
rect 22556 14660 22560 14716
rect 22496 14656 22560 14660
rect 28176 14716 28240 14720
rect 28176 14660 28180 14716
rect 28180 14660 28236 14716
rect 28236 14660 28240 14716
rect 28176 14656 28240 14660
rect 28256 14716 28320 14720
rect 28256 14660 28260 14716
rect 28260 14660 28316 14716
rect 28316 14660 28320 14716
rect 28256 14656 28320 14660
rect 28336 14716 28400 14720
rect 28336 14660 28340 14716
rect 28340 14660 28396 14716
rect 28396 14660 28400 14716
rect 28336 14656 28400 14660
rect 28416 14716 28480 14720
rect 28416 14660 28420 14716
rect 28420 14660 28476 14716
rect 28476 14660 28480 14716
rect 28416 14656 28480 14660
rect 28496 14716 28560 14720
rect 28496 14660 28500 14716
rect 28500 14660 28556 14716
rect 28556 14660 28560 14716
rect 28496 14656 28560 14660
rect 4916 14172 4980 14176
rect 4916 14116 4920 14172
rect 4920 14116 4976 14172
rect 4976 14116 4980 14172
rect 4916 14112 4980 14116
rect 4996 14172 5060 14176
rect 4996 14116 5000 14172
rect 5000 14116 5056 14172
rect 5056 14116 5060 14172
rect 4996 14112 5060 14116
rect 5076 14172 5140 14176
rect 5076 14116 5080 14172
rect 5080 14116 5136 14172
rect 5136 14116 5140 14172
rect 5076 14112 5140 14116
rect 5156 14172 5220 14176
rect 5156 14116 5160 14172
rect 5160 14116 5216 14172
rect 5216 14116 5220 14172
rect 5156 14112 5220 14116
rect 5236 14172 5300 14176
rect 5236 14116 5240 14172
rect 5240 14116 5296 14172
rect 5296 14116 5300 14172
rect 5236 14112 5300 14116
rect 10916 14172 10980 14176
rect 10916 14116 10920 14172
rect 10920 14116 10976 14172
rect 10976 14116 10980 14172
rect 10916 14112 10980 14116
rect 10996 14172 11060 14176
rect 10996 14116 11000 14172
rect 11000 14116 11056 14172
rect 11056 14116 11060 14172
rect 10996 14112 11060 14116
rect 11076 14172 11140 14176
rect 11076 14116 11080 14172
rect 11080 14116 11136 14172
rect 11136 14116 11140 14172
rect 11076 14112 11140 14116
rect 11156 14172 11220 14176
rect 11156 14116 11160 14172
rect 11160 14116 11216 14172
rect 11216 14116 11220 14172
rect 11156 14112 11220 14116
rect 11236 14172 11300 14176
rect 11236 14116 11240 14172
rect 11240 14116 11296 14172
rect 11296 14116 11300 14172
rect 11236 14112 11300 14116
rect 16916 14172 16980 14176
rect 16916 14116 16920 14172
rect 16920 14116 16976 14172
rect 16976 14116 16980 14172
rect 16916 14112 16980 14116
rect 16996 14172 17060 14176
rect 16996 14116 17000 14172
rect 17000 14116 17056 14172
rect 17056 14116 17060 14172
rect 16996 14112 17060 14116
rect 17076 14172 17140 14176
rect 17076 14116 17080 14172
rect 17080 14116 17136 14172
rect 17136 14116 17140 14172
rect 17076 14112 17140 14116
rect 17156 14172 17220 14176
rect 17156 14116 17160 14172
rect 17160 14116 17216 14172
rect 17216 14116 17220 14172
rect 17156 14112 17220 14116
rect 17236 14172 17300 14176
rect 17236 14116 17240 14172
rect 17240 14116 17296 14172
rect 17296 14116 17300 14172
rect 17236 14112 17300 14116
rect 22916 14172 22980 14176
rect 22916 14116 22920 14172
rect 22920 14116 22976 14172
rect 22976 14116 22980 14172
rect 22916 14112 22980 14116
rect 22996 14172 23060 14176
rect 22996 14116 23000 14172
rect 23000 14116 23056 14172
rect 23056 14116 23060 14172
rect 22996 14112 23060 14116
rect 23076 14172 23140 14176
rect 23076 14116 23080 14172
rect 23080 14116 23136 14172
rect 23136 14116 23140 14172
rect 23076 14112 23140 14116
rect 23156 14172 23220 14176
rect 23156 14116 23160 14172
rect 23160 14116 23216 14172
rect 23216 14116 23220 14172
rect 23156 14112 23220 14116
rect 23236 14172 23300 14176
rect 23236 14116 23240 14172
rect 23240 14116 23296 14172
rect 23296 14116 23300 14172
rect 23236 14112 23300 14116
rect 28916 14172 28980 14176
rect 28916 14116 28920 14172
rect 28920 14116 28976 14172
rect 28976 14116 28980 14172
rect 28916 14112 28980 14116
rect 28996 14172 29060 14176
rect 28996 14116 29000 14172
rect 29000 14116 29056 14172
rect 29056 14116 29060 14172
rect 28996 14112 29060 14116
rect 29076 14172 29140 14176
rect 29076 14116 29080 14172
rect 29080 14116 29136 14172
rect 29136 14116 29140 14172
rect 29076 14112 29140 14116
rect 29156 14172 29220 14176
rect 29156 14116 29160 14172
rect 29160 14116 29216 14172
rect 29216 14116 29220 14172
rect 29156 14112 29220 14116
rect 29236 14172 29300 14176
rect 29236 14116 29240 14172
rect 29240 14116 29296 14172
rect 29296 14116 29300 14172
rect 29236 14112 29300 14116
rect 4176 13628 4240 13632
rect 4176 13572 4180 13628
rect 4180 13572 4236 13628
rect 4236 13572 4240 13628
rect 4176 13568 4240 13572
rect 4256 13628 4320 13632
rect 4256 13572 4260 13628
rect 4260 13572 4316 13628
rect 4316 13572 4320 13628
rect 4256 13568 4320 13572
rect 4336 13628 4400 13632
rect 4336 13572 4340 13628
rect 4340 13572 4396 13628
rect 4396 13572 4400 13628
rect 4336 13568 4400 13572
rect 4416 13628 4480 13632
rect 4416 13572 4420 13628
rect 4420 13572 4476 13628
rect 4476 13572 4480 13628
rect 4416 13568 4480 13572
rect 4496 13628 4560 13632
rect 4496 13572 4500 13628
rect 4500 13572 4556 13628
rect 4556 13572 4560 13628
rect 4496 13568 4560 13572
rect 10176 13628 10240 13632
rect 10176 13572 10180 13628
rect 10180 13572 10236 13628
rect 10236 13572 10240 13628
rect 10176 13568 10240 13572
rect 10256 13628 10320 13632
rect 10256 13572 10260 13628
rect 10260 13572 10316 13628
rect 10316 13572 10320 13628
rect 10256 13568 10320 13572
rect 10336 13628 10400 13632
rect 10336 13572 10340 13628
rect 10340 13572 10396 13628
rect 10396 13572 10400 13628
rect 10336 13568 10400 13572
rect 10416 13628 10480 13632
rect 10416 13572 10420 13628
rect 10420 13572 10476 13628
rect 10476 13572 10480 13628
rect 10416 13568 10480 13572
rect 10496 13628 10560 13632
rect 10496 13572 10500 13628
rect 10500 13572 10556 13628
rect 10556 13572 10560 13628
rect 10496 13568 10560 13572
rect 16176 13628 16240 13632
rect 16176 13572 16180 13628
rect 16180 13572 16236 13628
rect 16236 13572 16240 13628
rect 16176 13568 16240 13572
rect 16256 13628 16320 13632
rect 16256 13572 16260 13628
rect 16260 13572 16316 13628
rect 16316 13572 16320 13628
rect 16256 13568 16320 13572
rect 16336 13628 16400 13632
rect 16336 13572 16340 13628
rect 16340 13572 16396 13628
rect 16396 13572 16400 13628
rect 16336 13568 16400 13572
rect 16416 13628 16480 13632
rect 16416 13572 16420 13628
rect 16420 13572 16476 13628
rect 16476 13572 16480 13628
rect 16416 13568 16480 13572
rect 16496 13628 16560 13632
rect 16496 13572 16500 13628
rect 16500 13572 16556 13628
rect 16556 13572 16560 13628
rect 16496 13568 16560 13572
rect 22176 13628 22240 13632
rect 22176 13572 22180 13628
rect 22180 13572 22236 13628
rect 22236 13572 22240 13628
rect 22176 13568 22240 13572
rect 22256 13628 22320 13632
rect 22256 13572 22260 13628
rect 22260 13572 22316 13628
rect 22316 13572 22320 13628
rect 22256 13568 22320 13572
rect 22336 13628 22400 13632
rect 22336 13572 22340 13628
rect 22340 13572 22396 13628
rect 22396 13572 22400 13628
rect 22336 13568 22400 13572
rect 22416 13628 22480 13632
rect 22416 13572 22420 13628
rect 22420 13572 22476 13628
rect 22476 13572 22480 13628
rect 22416 13568 22480 13572
rect 22496 13628 22560 13632
rect 22496 13572 22500 13628
rect 22500 13572 22556 13628
rect 22556 13572 22560 13628
rect 22496 13568 22560 13572
rect 28176 13628 28240 13632
rect 28176 13572 28180 13628
rect 28180 13572 28236 13628
rect 28236 13572 28240 13628
rect 28176 13568 28240 13572
rect 28256 13628 28320 13632
rect 28256 13572 28260 13628
rect 28260 13572 28316 13628
rect 28316 13572 28320 13628
rect 28256 13568 28320 13572
rect 28336 13628 28400 13632
rect 28336 13572 28340 13628
rect 28340 13572 28396 13628
rect 28396 13572 28400 13628
rect 28336 13568 28400 13572
rect 28416 13628 28480 13632
rect 28416 13572 28420 13628
rect 28420 13572 28476 13628
rect 28476 13572 28480 13628
rect 28416 13568 28480 13572
rect 28496 13628 28560 13632
rect 28496 13572 28500 13628
rect 28500 13572 28556 13628
rect 28556 13572 28560 13628
rect 28496 13568 28560 13572
rect 4916 13084 4980 13088
rect 4916 13028 4920 13084
rect 4920 13028 4976 13084
rect 4976 13028 4980 13084
rect 4916 13024 4980 13028
rect 4996 13084 5060 13088
rect 4996 13028 5000 13084
rect 5000 13028 5056 13084
rect 5056 13028 5060 13084
rect 4996 13024 5060 13028
rect 5076 13084 5140 13088
rect 5076 13028 5080 13084
rect 5080 13028 5136 13084
rect 5136 13028 5140 13084
rect 5076 13024 5140 13028
rect 5156 13084 5220 13088
rect 5156 13028 5160 13084
rect 5160 13028 5216 13084
rect 5216 13028 5220 13084
rect 5156 13024 5220 13028
rect 5236 13084 5300 13088
rect 5236 13028 5240 13084
rect 5240 13028 5296 13084
rect 5296 13028 5300 13084
rect 5236 13024 5300 13028
rect 10916 13084 10980 13088
rect 10916 13028 10920 13084
rect 10920 13028 10976 13084
rect 10976 13028 10980 13084
rect 10916 13024 10980 13028
rect 10996 13084 11060 13088
rect 10996 13028 11000 13084
rect 11000 13028 11056 13084
rect 11056 13028 11060 13084
rect 10996 13024 11060 13028
rect 11076 13084 11140 13088
rect 11076 13028 11080 13084
rect 11080 13028 11136 13084
rect 11136 13028 11140 13084
rect 11076 13024 11140 13028
rect 11156 13084 11220 13088
rect 11156 13028 11160 13084
rect 11160 13028 11216 13084
rect 11216 13028 11220 13084
rect 11156 13024 11220 13028
rect 11236 13084 11300 13088
rect 11236 13028 11240 13084
rect 11240 13028 11296 13084
rect 11296 13028 11300 13084
rect 11236 13024 11300 13028
rect 16916 13084 16980 13088
rect 16916 13028 16920 13084
rect 16920 13028 16976 13084
rect 16976 13028 16980 13084
rect 16916 13024 16980 13028
rect 16996 13084 17060 13088
rect 16996 13028 17000 13084
rect 17000 13028 17056 13084
rect 17056 13028 17060 13084
rect 16996 13024 17060 13028
rect 17076 13084 17140 13088
rect 17076 13028 17080 13084
rect 17080 13028 17136 13084
rect 17136 13028 17140 13084
rect 17076 13024 17140 13028
rect 17156 13084 17220 13088
rect 17156 13028 17160 13084
rect 17160 13028 17216 13084
rect 17216 13028 17220 13084
rect 17156 13024 17220 13028
rect 17236 13084 17300 13088
rect 17236 13028 17240 13084
rect 17240 13028 17296 13084
rect 17296 13028 17300 13084
rect 17236 13024 17300 13028
rect 22916 13084 22980 13088
rect 22916 13028 22920 13084
rect 22920 13028 22976 13084
rect 22976 13028 22980 13084
rect 22916 13024 22980 13028
rect 22996 13084 23060 13088
rect 22996 13028 23000 13084
rect 23000 13028 23056 13084
rect 23056 13028 23060 13084
rect 22996 13024 23060 13028
rect 23076 13084 23140 13088
rect 23076 13028 23080 13084
rect 23080 13028 23136 13084
rect 23136 13028 23140 13084
rect 23076 13024 23140 13028
rect 23156 13084 23220 13088
rect 23156 13028 23160 13084
rect 23160 13028 23216 13084
rect 23216 13028 23220 13084
rect 23156 13024 23220 13028
rect 23236 13084 23300 13088
rect 23236 13028 23240 13084
rect 23240 13028 23296 13084
rect 23296 13028 23300 13084
rect 23236 13024 23300 13028
rect 28916 13084 28980 13088
rect 28916 13028 28920 13084
rect 28920 13028 28976 13084
rect 28976 13028 28980 13084
rect 28916 13024 28980 13028
rect 28996 13084 29060 13088
rect 28996 13028 29000 13084
rect 29000 13028 29056 13084
rect 29056 13028 29060 13084
rect 28996 13024 29060 13028
rect 29076 13084 29140 13088
rect 29076 13028 29080 13084
rect 29080 13028 29136 13084
rect 29136 13028 29140 13084
rect 29076 13024 29140 13028
rect 29156 13084 29220 13088
rect 29156 13028 29160 13084
rect 29160 13028 29216 13084
rect 29216 13028 29220 13084
rect 29156 13024 29220 13028
rect 29236 13084 29300 13088
rect 29236 13028 29240 13084
rect 29240 13028 29296 13084
rect 29296 13028 29300 13084
rect 29236 13024 29300 13028
rect 15332 12820 15396 12884
rect 4176 12540 4240 12544
rect 4176 12484 4180 12540
rect 4180 12484 4236 12540
rect 4236 12484 4240 12540
rect 4176 12480 4240 12484
rect 4256 12540 4320 12544
rect 4256 12484 4260 12540
rect 4260 12484 4316 12540
rect 4316 12484 4320 12540
rect 4256 12480 4320 12484
rect 4336 12540 4400 12544
rect 4336 12484 4340 12540
rect 4340 12484 4396 12540
rect 4396 12484 4400 12540
rect 4336 12480 4400 12484
rect 4416 12540 4480 12544
rect 4416 12484 4420 12540
rect 4420 12484 4476 12540
rect 4476 12484 4480 12540
rect 4416 12480 4480 12484
rect 4496 12540 4560 12544
rect 4496 12484 4500 12540
rect 4500 12484 4556 12540
rect 4556 12484 4560 12540
rect 4496 12480 4560 12484
rect 10176 12540 10240 12544
rect 10176 12484 10180 12540
rect 10180 12484 10236 12540
rect 10236 12484 10240 12540
rect 10176 12480 10240 12484
rect 10256 12540 10320 12544
rect 10256 12484 10260 12540
rect 10260 12484 10316 12540
rect 10316 12484 10320 12540
rect 10256 12480 10320 12484
rect 10336 12540 10400 12544
rect 10336 12484 10340 12540
rect 10340 12484 10396 12540
rect 10396 12484 10400 12540
rect 10336 12480 10400 12484
rect 10416 12540 10480 12544
rect 10416 12484 10420 12540
rect 10420 12484 10476 12540
rect 10476 12484 10480 12540
rect 10416 12480 10480 12484
rect 10496 12540 10560 12544
rect 10496 12484 10500 12540
rect 10500 12484 10556 12540
rect 10556 12484 10560 12540
rect 10496 12480 10560 12484
rect 16176 12540 16240 12544
rect 16176 12484 16180 12540
rect 16180 12484 16236 12540
rect 16236 12484 16240 12540
rect 16176 12480 16240 12484
rect 16256 12540 16320 12544
rect 16256 12484 16260 12540
rect 16260 12484 16316 12540
rect 16316 12484 16320 12540
rect 16256 12480 16320 12484
rect 16336 12540 16400 12544
rect 16336 12484 16340 12540
rect 16340 12484 16396 12540
rect 16396 12484 16400 12540
rect 16336 12480 16400 12484
rect 16416 12540 16480 12544
rect 16416 12484 16420 12540
rect 16420 12484 16476 12540
rect 16476 12484 16480 12540
rect 16416 12480 16480 12484
rect 16496 12540 16560 12544
rect 16496 12484 16500 12540
rect 16500 12484 16556 12540
rect 16556 12484 16560 12540
rect 16496 12480 16560 12484
rect 22176 12540 22240 12544
rect 22176 12484 22180 12540
rect 22180 12484 22236 12540
rect 22236 12484 22240 12540
rect 22176 12480 22240 12484
rect 22256 12540 22320 12544
rect 22256 12484 22260 12540
rect 22260 12484 22316 12540
rect 22316 12484 22320 12540
rect 22256 12480 22320 12484
rect 22336 12540 22400 12544
rect 22336 12484 22340 12540
rect 22340 12484 22396 12540
rect 22396 12484 22400 12540
rect 22336 12480 22400 12484
rect 22416 12540 22480 12544
rect 22416 12484 22420 12540
rect 22420 12484 22476 12540
rect 22476 12484 22480 12540
rect 22416 12480 22480 12484
rect 22496 12540 22560 12544
rect 22496 12484 22500 12540
rect 22500 12484 22556 12540
rect 22556 12484 22560 12540
rect 22496 12480 22560 12484
rect 28176 12540 28240 12544
rect 28176 12484 28180 12540
rect 28180 12484 28236 12540
rect 28236 12484 28240 12540
rect 28176 12480 28240 12484
rect 28256 12540 28320 12544
rect 28256 12484 28260 12540
rect 28260 12484 28316 12540
rect 28316 12484 28320 12540
rect 28256 12480 28320 12484
rect 28336 12540 28400 12544
rect 28336 12484 28340 12540
rect 28340 12484 28396 12540
rect 28396 12484 28400 12540
rect 28336 12480 28400 12484
rect 28416 12540 28480 12544
rect 28416 12484 28420 12540
rect 28420 12484 28476 12540
rect 28476 12484 28480 12540
rect 28416 12480 28480 12484
rect 28496 12540 28560 12544
rect 28496 12484 28500 12540
rect 28500 12484 28556 12540
rect 28556 12484 28560 12540
rect 28496 12480 28560 12484
rect 4916 11996 4980 12000
rect 4916 11940 4920 11996
rect 4920 11940 4976 11996
rect 4976 11940 4980 11996
rect 4916 11936 4980 11940
rect 4996 11996 5060 12000
rect 4996 11940 5000 11996
rect 5000 11940 5056 11996
rect 5056 11940 5060 11996
rect 4996 11936 5060 11940
rect 5076 11996 5140 12000
rect 5076 11940 5080 11996
rect 5080 11940 5136 11996
rect 5136 11940 5140 11996
rect 5076 11936 5140 11940
rect 5156 11996 5220 12000
rect 5156 11940 5160 11996
rect 5160 11940 5216 11996
rect 5216 11940 5220 11996
rect 5156 11936 5220 11940
rect 5236 11996 5300 12000
rect 5236 11940 5240 11996
rect 5240 11940 5296 11996
rect 5296 11940 5300 11996
rect 5236 11936 5300 11940
rect 10916 11996 10980 12000
rect 10916 11940 10920 11996
rect 10920 11940 10976 11996
rect 10976 11940 10980 11996
rect 10916 11936 10980 11940
rect 10996 11996 11060 12000
rect 10996 11940 11000 11996
rect 11000 11940 11056 11996
rect 11056 11940 11060 11996
rect 10996 11936 11060 11940
rect 11076 11996 11140 12000
rect 11076 11940 11080 11996
rect 11080 11940 11136 11996
rect 11136 11940 11140 11996
rect 11076 11936 11140 11940
rect 11156 11996 11220 12000
rect 11156 11940 11160 11996
rect 11160 11940 11216 11996
rect 11216 11940 11220 11996
rect 11156 11936 11220 11940
rect 11236 11996 11300 12000
rect 11236 11940 11240 11996
rect 11240 11940 11296 11996
rect 11296 11940 11300 11996
rect 11236 11936 11300 11940
rect 16916 11996 16980 12000
rect 16916 11940 16920 11996
rect 16920 11940 16976 11996
rect 16976 11940 16980 11996
rect 16916 11936 16980 11940
rect 16996 11996 17060 12000
rect 16996 11940 17000 11996
rect 17000 11940 17056 11996
rect 17056 11940 17060 11996
rect 16996 11936 17060 11940
rect 17076 11996 17140 12000
rect 17076 11940 17080 11996
rect 17080 11940 17136 11996
rect 17136 11940 17140 11996
rect 17076 11936 17140 11940
rect 17156 11996 17220 12000
rect 17156 11940 17160 11996
rect 17160 11940 17216 11996
rect 17216 11940 17220 11996
rect 17156 11936 17220 11940
rect 17236 11996 17300 12000
rect 17236 11940 17240 11996
rect 17240 11940 17296 11996
rect 17296 11940 17300 11996
rect 17236 11936 17300 11940
rect 22916 11996 22980 12000
rect 22916 11940 22920 11996
rect 22920 11940 22976 11996
rect 22976 11940 22980 11996
rect 22916 11936 22980 11940
rect 22996 11996 23060 12000
rect 22996 11940 23000 11996
rect 23000 11940 23056 11996
rect 23056 11940 23060 11996
rect 22996 11936 23060 11940
rect 23076 11996 23140 12000
rect 23076 11940 23080 11996
rect 23080 11940 23136 11996
rect 23136 11940 23140 11996
rect 23076 11936 23140 11940
rect 23156 11996 23220 12000
rect 23156 11940 23160 11996
rect 23160 11940 23216 11996
rect 23216 11940 23220 11996
rect 23156 11936 23220 11940
rect 23236 11996 23300 12000
rect 23236 11940 23240 11996
rect 23240 11940 23296 11996
rect 23296 11940 23300 11996
rect 23236 11936 23300 11940
rect 28916 11996 28980 12000
rect 28916 11940 28920 11996
rect 28920 11940 28976 11996
rect 28976 11940 28980 11996
rect 28916 11936 28980 11940
rect 28996 11996 29060 12000
rect 28996 11940 29000 11996
rect 29000 11940 29056 11996
rect 29056 11940 29060 11996
rect 28996 11936 29060 11940
rect 29076 11996 29140 12000
rect 29076 11940 29080 11996
rect 29080 11940 29136 11996
rect 29136 11940 29140 11996
rect 29076 11936 29140 11940
rect 29156 11996 29220 12000
rect 29156 11940 29160 11996
rect 29160 11940 29216 11996
rect 29216 11940 29220 11996
rect 29156 11936 29220 11940
rect 29236 11996 29300 12000
rect 29236 11940 29240 11996
rect 29240 11940 29296 11996
rect 29296 11940 29300 11996
rect 29236 11936 29300 11940
rect 4176 11452 4240 11456
rect 4176 11396 4180 11452
rect 4180 11396 4236 11452
rect 4236 11396 4240 11452
rect 4176 11392 4240 11396
rect 4256 11452 4320 11456
rect 4256 11396 4260 11452
rect 4260 11396 4316 11452
rect 4316 11396 4320 11452
rect 4256 11392 4320 11396
rect 4336 11452 4400 11456
rect 4336 11396 4340 11452
rect 4340 11396 4396 11452
rect 4396 11396 4400 11452
rect 4336 11392 4400 11396
rect 4416 11452 4480 11456
rect 4416 11396 4420 11452
rect 4420 11396 4476 11452
rect 4476 11396 4480 11452
rect 4416 11392 4480 11396
rect 4496 11452 4560 11456
rect 4496 11396 4500 11452
rect 4500 11396 4556 11452
rect 4556 11396 4560 11452
rect 4496 11392 4560 11396
rect 10176 11452 10240 11456
rect 10176 11396 10180 11452
rect 10180 11396 10236 11452
rect 10236 11396 10240 11452
rect 10176 11392 10240 11396
rect 10256 11452 10320 11456
rect 10256 11396 10260 11452
rect 10260 11396 10316 11452
rect 10316 11396 10320 11452
rect 10256 11392 10320 11396
rect 10336 11452 10400 11456
rect 10336 11396 10340 11452
rect 10340 11396 10396 11452
rect 10396 11396 10400 11452
rect 10336 11392 10400 11396
rect 10416 11452 10480 11456
rect 10416 11396 10420 11452
rect 10420 11396 10476 11452
rect 10476 11396 10480 11452
rect 10416 11392 10480 11396
rect 10496 11452 10560 11456
rect 10496 11396 10500 11452
rect 10500 11396 10556 11452
rect 10556 11396 10560 11452
rect 10496 11392 10560 11396
rect 16176 11452 16240 11456
rect 16176 11396 16180 11452
rect 16180 11396 16236 11452
rect 16236 11396 16240 11452
rect 16176 11392 16240 11396
rect 16256 11452 16320 11456
rect 16256 11396 16260 11452
rect 16260 11396 16316 11452
rect 16316 11396 16320 11452
rect 16256 11392 16320 11396
rect 16336 11452 16400 11456
rect 16336 11396 16340 11452
rect 16340 11396 16396 11452
rect 16396 11396 16400 11452
rect 16336 11392 16400 11396
rect 16416 11452 16480 11456
rect 16416 11396 16420 11452
rect 16420 11396 16476 11452
rect 16476 11396 16480 11452
rect 16416 11392 16480 11396
rect 16496 11452 16560 11456
rect 16496 11396 16500 11452
rect 16500 11396 16556 11452
rect 16556 11396 16560 11452
rect 16496 11392 16560 11396
rect 22176 11452 22240 11456
rect 22176 11396 22180 11452
rect 22180 11396 22236 11452
rect 22236 11396 22240 11452
rect 22176 11392 22240 11396
rect 22256 11452 22320 11456
rect 22256 11396 22260 11452
rect 22260 11396 22316 11452
rect 22316 11396 22320 11452
rect 22256 11392 22320 11396
rect 22336 11452 22400 11456
rect 22336 11396 22340 11452
rect 22340 11396 22396 11452
rect 22396 11396 22400 11452
rect 22336 11392 22400 11396
rect 22416 11452 22480 11456
rect 22416 11396 22420 11452
rect 22420 11396 22476 11452
rect 22476 11396 22480 11452
rect 22416 11392 22480 11396
rect 22496 11452 22560 11456
rect 22496 11396 22500 11452
rect 22500 11396 22556 11452
rect 22556 11396 22560 11452
rect 22496 11392 22560 11396
rect 28176 11452 28240 11456
rect 28176 11396 28180 11452
rect 28180 11396 28236 11452
rect 28236 11396 28240 11452
rect 28176 11392 28240 11396
rect 28256 11452 28320 11456
rect 28256 11396 28260 11452
rect 28260 11396 28316 11452
rect 28316 11396 28320 11452
rect 28256 11392 28320 11396
rect 28336 11452 28400 11456
rect 28336 11396 28340 11452
rect 28340 11396 28396 11452
rect 28396 11396 28400 11452
rect 28336 11392 28400 11396
rect 28416 11452 28480 11456
rect 28416 11396 28420 11452
rect 28420 11396 28476 11452
rect 28476 11396 28480 11452
rect 28416 11392 28480 11396
rect 28496 11452 28560 11456
rect 28496 11396 28500 11452
rect 28500 11396 28556 11452
rect 28556 11396 28560 11452
rect 28496 11392 28560 11396
rect 15332 11112 15396 11116
rect 15332 11056 15382 11112
rect 15382 11056 15396 11112
rect 15332 11052 15396 11056
rect 4916 10908 4980 10912
rect 4916 10852 4920 10908
rect 4920 10852 4976 10908
rect 4976 10852 4980 10908
rect 4916 10848 4980 10852
rect 4996 10908 5060 10912
rect 4996 10852 5000 10908
rect 5000 10852 5056 10908
rect 5056 10852 5060 10908
rect 4996 10848 5060 10852
rect 5076 10908 5140 10912
rect 5076 10852 5080 10908
rect 5080 10852 5136 10908
rect 5136 10852 5140 10908
rect 5076 10848 5140 10852
rect 5156 10908 5220 10912
rect 5156 10852 5160 10908
rect 5160 10852 5216 10908
rect 5216 10852 5220 10908
rect 5156 10848 5220 10852
rect 5236 10908 5300 10912
rect 5236 10852 5240 10908
rect 5240 10852 5296 10908
rect 5296 10852 5300 10908
rect 5236 10848 5300 10852
rect 10916 10908 10980 10912
rect 10916 10852 10920 10908
rect 10920 10852 10976 10908
rect 10976 10852 10980 10908
rect 10916 10848 10980 10852
rect 10996 10908 11060 10912
rect 10996 10852 11000 10908
rect 11000 10852 11056 10908
rect 11056 10852 11060 10908
rect 10996 10848 11060 10852
rect 11076 10908 11140 10912
rect 11076 10852 11080 10908
rect 11080 10852 11136 10908
rect 11136 10852 11140 10908
rect 11076 10848 11140 10852
rect 11156 10908 11220 10912
rect 11156 10852 11160 10908
rect 11160 10852 11216 10908
rect 11216 10852 11220 10908
rect 11156 10848 11220 10852
rect 11236 10908 11300 10912
rect 11236 10852 11240 10908
rect 11240 10852 11296 10908
rect 11296 10852 11300 10908
rect 11236 10848 11300 10852
rect 16916 10908 16980 10912
rect 16916 10852 16920 10908
rect 16920 10852 16976 10908
rect 16976 10852 16980 10908
rect 16916 10848 16980 10852
rect 16996 10908 17060 10912
rect 16996 10852 17000 10908
rect 17000 10852 17056 10908
rect 17056 10852 17060 10908
rect 16996 10848 17060 10852
rect 17076 10908 17140 10912
rect 17076 10852 17080 10908
rect 17080 10852 17136 10908
rect 17136 10852 17140 10908
rect 17076 10848 17140 10852
rect 17156 10908 17220 10912
rect 17156 10852 17160 10908
rect 17160 10852 17216 10908
rect 17216 10852 17220 10908
rect 17156 10848 17220 10852
rect 17236 10908 17300 10912
rect 17236 10852 17240 10908
rect 17240 10852 17296 10908
rect 17296 10852 17300 10908
rect 17236 10848 17300 10852
rect 22916 10908 22980 10912
rect 22916 10852 22920 10908
rect 22920 10852 22976 10908
rect 22976 10852 22980 10908
rect 22916 10848 22980 10852
rect 22996 10908 23060 10912
rect 22996 10852 23000 10908
rect 23000 10852 23056 10908
rect 23056 10852 23060 10908
rect 22996 10848 23060 10852
rect 23076 10908 23140 10912
rect 23076 10852 23080 10908
rect 23080 10852 23136 10908
rect 23136 10852 23140 10908
rect 23076 10848 23140 10852
rect 23156 10908 23220 10912
rect 23156 10852 23160 10908
rect 23160 10852 23216 10908
rect 23216 10852 23220 10908
rect 23156 10848 23220 10852
rect 23236 10908 23300 10912
rect 23236 10852 23240 10908
rect 23240 10852 23296 10908
rect 23296 10852 23300 10908
rect 23236 10848 23300 10852
rect 28916 10908 28980 10912
rect 28916 10852 28920 10908
rect 28920 10852 28976 10908
rect 28976 10852 28980 10908
rect 28916 10848 28980 10852
rect 28996 10908 29060 10912
rect 28996 10852 29000 10908
rect 29000 10852 29056 10908
rect 29056 10852 29060 10908
rect 28996 10848 29060 10852
rect 29076 10908 29140 10912
rect 29076 10852 29080 10908
rect 29080 10852 29136 10908
rect 29136 10852 29140 10908
rect 29076 10848 29140 10852
rect 29156 10908 29220 10912
rect 29156 10852 29160 10908
rect 29160 10852 29216 10908
rect 29216 10852 29220 10908
rect 29156 10848 29220 10852
rect 29236 10908 29300 10912
rect 29236 10852 29240 10908
rect 29240 10852 29296 10908
rect 29296 10852 29300 10908
rect 29236 10848 29300 10852
rect 4176 10364 4240 10368
rect 4176 10308 4180 10364
rect 4180 10308 4236 10364
rect 4236 10308 4240 10364
rect 4176 10304 4240 10308
rect 4256 10364 4320 10368
rect 4256 10308 4260 10364
rect 4260 10308 4316 10364
rect 4316 10308 4320 10364
rect 4256 10304 4320 10308
rect 4336 10364 4400 10368
rect 4336 10308 4340 10364
rect 4340 10308 4396 10364
rect 4396 10308 4400 10364
rect 4336 10304 4400 10308
rect 4416 10364 4480 10368
rect 4416 10308 4420 10364
rect 4420 10308 4476 10364
rect 4476 10308 4480 10364
rect 4416 10304 4480 10308
rect 4496 10364 4560 10368
rect 4496 10308 4500 10364
rect 4500 10308 4556 10364
rect 4556 10308 4560 10364
rect 4496 10304 4560 10308
rect 10176 10364 10240 10368
rect 10176 10308 10180 10364
rect 10180 10308 10236 10364
rect 10236 10308 10240 10364
rect 10176 10304 10240 10308
rect 10256 10364 10320 10368
rect 10256 10308 10260 10364
rect 10260 10308 10316 10364
rect 10316 10308 10320 10364
rect 10256 10304 10320 10308
rect 10336 10364 10400 10368
rect 10336 10308 10340 10364
rect 10340 10308 10396 10364
rect 10396 10308 10400 10364
rect 10336 10304 10400 10308
rect 10416 10364 10480 10368
rect 10416 10308 10420 10364
rect 10420 10308 10476 10364
rect 10476 10308 10480 10364
rect 10416 10304 10480 10308
rect 10496 10364 10560 10368
rect 10496 10308 10500 10364
rect 10500 10308 10556 10364
rect 10556 10308 10560 10364
rect 10496 10304 10560 10308
rect 16176 10364 16240 10368
rect 16176 10308 16180 10364
rect 16180 10308 16236 10364
rect 16236 10308 16240 10364
rect 16176 10304 16240 10308
rect 16256 10364 16320 10368
rect 16256 10308 16260 10364
rect 16260 10308 16316 10364
rect 16316 10308 16320 10364
rect 16256 10304 16320 10308
rect 16336 10364 16400 10368
rect 16336 10308 16340 10364
rect 16340 10308 16396 10364
rect 16396 10308 16400 10364
rect 16336 10304 16400 10308
rect 16416 10364 16480 10368
rect 16416 10308 16420 10364
rect 16420 10308 16476 10364
rect 16476 10308 16480 10364
rect 16416 10304 16480 10308
rect 16496 10364 16560 10368
rect 16496 10308 16500 10364
rect 16500 10308 16556 10364
rect 16556 10308 16560 10364
rect 16496 10304 16560 10308
rect 22176 10364 22240 10368
rect 22176 10308 22180 10364
rect 22180 10308 22236 10364
rect 22236 10308 22240 10364
rect 22176 10304 22240 10308
rect 22256 10364 22320 10368
rect 22256 10308 22260 10364
rect 22260 10308 22316 10364
rect 22316 10308 22320 10364
rect 22256 10304 22320 10308
rect 22336 10364 22400 10368
rect 22336 10308 22340 10364
rect 22340 10308 22396 10364
rect 22396 10308 22400 10364
rect 22336 10304 22400 10308
rect 22416 10364 22480 10368
rect 22416 10308 22420 10364
rect 22420 10308 22476 10364
rect 22476 10308 22480 10364
rect 22416 10304 22480 10308
rect 22496 10364 22560 10368
rect 22496 10308 22500 10364
rect 22500 10308 22556 10364
rect 22556 10308 22560 10364
rect 22496 10304 22560 10308
rect 28176 10364 28240 10368
rect 28176 10308 28180 10364
rect 28180 10308 28236 10364
rect 28236 10308 28240 10364
rect 28176 10304 28240 10308
rect 28256 10364 28320 10368
rect 28256 10308 28260 10364
rect 28260 10308 28316 10364
rect 28316 10308 28320 10364
rect 28256 10304 28320 10308
rect 28336 10364 28400 10368
rect 28336 10308 28340 10364
rect 28340 10308 28396 10364
rect 28396 10308 28400 10364
rect 28336 10304 28400 10308
rect 28416 10364 28480 10368
rect 28416 10308 28420 10364
rect 28420 10308 28476 10364
rect 28476 10308 28480 10364
rect 28416 10304 28480 10308
rect 28496 10364 28560 10368
rect 28496 10308 28500 10364
rect 28500 10308 28556 10364
rect 28556 10308 28560 10364
rect 28496 10304 28560 10308
rect 4916 9820 4980 9824
rect 4916 9764 4920 9820
rect 4920 9764 4976 9820
rect 4976 9764 4980 9820
rect 4916 9760 4980 9764
rect 4996 9820 5060 9824
rect 4996 9764 5000 9820
rect 5000 9764 5056 9820
rect 5056 9764 5060 9820
rect 4996 9760 5060 9764
rect 5076 9820 5140 9824
rect 5076 9764 5080 9820
rect 5080 9764 5136 9820
rect 5136 9764 5140 9820
rect 5076 9760 5140 9764
rect 5156 9820 5220 9824
rect 5156 9764 5160 9820
rect 5160 9764 5216 9820
rect 5216 9764 5220 9820
rect 5156 9760 5220 9764
rect 5236 9820 5300 9824
rect 5236 9764 5240 9820
rect 5240 9764 5296 9820
rect 5296 9764 5300 9820
rect 5236 9760 5300 9764
rect 10916 9820 10980 9824
rect 10916 9764 10920 9820
rect 10920 9764 10976 9820
rect 10976 9764 10980 9820
rect 10916 9760 10980 9764
rect 10996 9820 11060 9824
rect 10996 9764 11000 9820
rect 11000 9764 11056 9820
rect 11056 9764 11060 9820
rect 10996 9760 11060 9764
rect 11076 9820 11140 9824
rect 11076 9764 11080 9820
rect 11080 9764 11136 9820
rect 11136 9764 11140 9820
rect 11076 9760 11140 9764
rect 11156 9820 11220 9824
rect 11156 9764 11160 9820
rect 11160 9764 11216 9820
rect 11216 9764 11220 9820
rect 11156 9760 11220 9764
rect 11236 9820 11300 9824
rect 11236 9764 11240 9820
rect 11240 9764 11296 9820
rect 11296 9764 11300 9820
rect 11236 9760 11300 9764
rect 16916 9820 16980 9824
rect 16916 9764 16920 9820
rect 16920 9764 16976 9820
rect 16976 9764 16980 9820
rect 16916 9760 16980 9764
rect 16996 9820 17060 9824
rect 16996 9764 17000 9820
rect 17000 9764 17056 9820
rect 17056 9764 17060 9820
rect 16996 9760 17060 9764
rect 17076 9820 17140 9824
rect 17076 9764 17080 9820
rect 17080 9764 17136 9820
rect 17136 9764 17140 9820
rect 17076 9760 17140 9764
rect 17156 9820 17220 9824
rect 17156 9764 17160 9820
rect 17160 9764 17216 9820
rect 17216 9764 17220 9820
rect 17156 9760 17220 9764
rect 17236 9820 17300 9824
rect 17236 9764 17240 9820
rect 17240 9764 17296 9820
rect 17296 9764 17300 9820
rect 17236 9760 17300 9764
rect 22916 9820 22980 9824
rect 22916 9764 22920 9820
rect 22920 9764 22976 9820
rect 22976 9764 22980 9820
rect 22916 9760 22980 9764
rect 22996 9820 23060 9824
rect 22996 9764 23000 9820
rect 23000 9764 23056 9820
rect 23056 9764 23060 9820
rect 22996 9760 23060 9764
rect 23076 9820 23140 9824
rect 23076 9764 23080 9820
rect 23080 9764 23136 9820
rect 23136 9764 23140 9820
rect 23076 9760 23140 9764
rect 23156 9820 23220 9824
rect 23156 9764 23160 9820
rect 23160 9764 23216 9820
rect 23216 9764 23220 9820
rect 23156 9760 23220 9764
rect 23236 9820 23300 9824
rect 23236 9764 23240 9820
rect 23240 9764 23296 9820
rect 23296 9764 23300 9820
rect 23236 9760 23300 9764
rect 28916 9820 28980 9824
rect 28916 9764 28920 9820
rect 28920 9764 28976 9820
rect 28976 9764 28980 9820
rect 28916 9760 28980 9764
rect 28996 9820 29060 9824
rect 28996 9764 29000 9820
rect 29000 9764 29056 9820
rect 29056 9764 29060 9820
rect 28996 9760 29060 9764
rect 29076 9820 29140 9824
rect 29076 9764 29080 9820
rect 29080 9764 29136 9820
rect 29136 9764 29140 9820
rect 29076 9760 29140 9764
rect 29156 9820 29220 9824
rect 29156 9764 29160 9820
rect 29160 9764 29216 9820
rect 29216 9764 29220 9820
rect 29156 9760 29220 9764
rect 29236 9820 29300 9824
rect 29236 9764 29240 9820
rect 29240 9764 29296 9820
rect 29296 9764 29300 9820
rect 29236 9760 29300 9764
rect 4176 9276 4240 9280
rect 4176 9220 4180 9276
rect 4180 9220 4236 9276
rect 4236 9220 4240 9276
rect 4176 9216 4240 9220
rect 4256 9276 4320 9280
rect 4256 9220 4260 9276
rect 4260 9220 4316 9276
rect 4316 9220 4320 9276
rect 4256 9216 4320 9220
rect 4336 9276 4400 9280
rect 4336 9220 4340 9276
rect 4340 9220 4396 9276
rect 4396 9220 4400 9276
rect 4336 9216 4400 9220
rect 4416 9276 4480 9280
rect 4416 9220 4420 9276
rect 4420 9220 4476 9276
rect 4476 9220 4480 9276
rect 4416 9216 4480 9220
rect 4496 9276 4560 9280
rect 4496 9220 4500 9276
rect 4500 9220 4556 9276
rect 4556 9220 4560 9276
rect 4496 9216 4560 9220
rect 10176 9276 10240 9280
rect 10176 9220 10180 9276
rect 10180 9220 10236 9276
rect 10236 9220 10240 9276
rect 10176 9216 10240 9220
rect 10256 9276 10320 9280
rect 10256 9220 10260 9276
rect 10260 9220 10316 9276
rect 10316 9220 10320 9276
rect 10256 9216 10320 9220
rect 10336 9276 10400 9280
rect 10336 9220 10340 9276
rect 10340 9220 10396 9276
rect 10396 9220 10400 9276
rect 10336 9216 10400 9220
rect 10416 9276 10480 9280
rect 10416 9220 10420 9276
rect 10420 9220 10476 9276
rect 10476 9220 10480 9276
rect 10416 9216 10480 9220
rect 10496 9276 10560 9280
rect 10496 9220 10500 9276
rect 10500 9220 10556 9276
rect 10556 9220 10560 9276
rect 10496 9216 10560 9220
rect 16176 9276 16240 9280
rect 16176 9220 16180 9276
rect 16180 9220 16236 9276
rect 16236 9220 16240 9276
rect 16176 9216 16240 9220
rect 16256 9276 16320 9280
rect 16256 9220 16260 9276
rect 16260 9220 16316 9276
rect 16316 9220 16320 9276
rect 16256 9216 16320 9220
rect 16336 9276 16400 9280
rect 16336 9220 16340 9276
rect 16340 9220 16396 9276
rect 16396 9220 16400 9276
rect 16336 9216 16400 9220
rect 16416 9276 16480 9280
rect 16416 9220 16420 9276
rect 16420 9220 16476 9276
rect 16476 9220 16480 9276
rect 16416 9216 16480 9220
rect 16496 9276 16560 9280
rect 16496 9220 16500 9276
rect 16500 9220 16556 9276
rect 16556 9220 16560 9276
rect 16496 9216 16560 9220
rect 22176 9276 22240 9280
rect 22176 9220 22180 9276
rect 22180 9220 22236 9276
rect 22236 9220 22240 9276
rect 22176 9216 22240 9220
rect 22256 9276 22320 9280
rect 22256 9220 22260 9276
rect 22260 9220 22316 9276
rect 22316 9220 22320 9276
rect 22256 9216 22320 9220
rect 22336 9276 22400 9280
rect 22336 9220 22340 9276
rect 22340 9220 22396 9276
rect 22396 9220 22400 9276
rect 22336 9216 22400 9220
rect 22416 9276 22480 9280
rect 22416 9220 22420 9276
rect 22420 9220 22476 9276
rect 22476 9220 22480 9276
rect 22416 9216 22480 9220
rect 22496 9276 22560 9280
rect 22496 9220 22500 9276
rect 22500 9220 22556 9276
rect 22556 9220 22560 9276
rect 22496 9216 22560 9220
rect 28176 9276 28240 9280
rect 28176 9220 28180 9276
rect 28180 9220 28236 9276
rect 28236 9220 28240 9276
rect 28176 9216 28240 9220
rect 28256 9276 28320 9280
rect 28256 9220 28260 9276
rect 28260 9220 28316 9276
rect 28316 9220 28320 9276
rect 28256 9216 28320 9220
rect 28336 9276 28400 9280
rect 28336 9220 28340 9276
rect 28340 9220 28396 9276
rect 28396 9220 28400 9276
rect 28336 9216 28400 9220
rect 28416 9276 28480 9280
rect 28416 9220 28420 9276
rect 28420 9220 28476 9276
rect 28476 9220 28480 9276
rect 28416 9216 28480 9220
rect 28496 9276 28560 9280
rect 28496 9220 28500 9276
rect 28500 9220 28556 9276
rect 28556 9220 28560 9276
rect 28496 9216 28560 9220
rect 18644 8740 18708 8804
rect 4916 8732 4980 8736
rect 4916 8676 4920 8732
rect 4920 8676 4976 8732
rect 4976 8676 4980 8732
rect 4916 8672 4980 8676
rect 4996 8732 5060 8736
rect 4996 8676 5000 8732
rect 5000 8676 5056 8732
rect 5056 8676 5060 8732
rect 4996 8672 5060 8676
rect 5076 8732 5140 8736
rect 5076 8676 5080 8732
rect 5080 8676 5136 8732
rect 5136 8676 5140 8732
rect 5076 8672 5140 8676
rect 5156 8732 5220 8736
rect 5156 8676 5160 8732
rect 5160 8676 5216 8732
rect 5216 8676 5220 8732
rect 5156 8672 5220 8676
rect 5236 8732 5300 8736
rect 5236 8676 5240 8732
rect 5240 8676 5296 8732
rect 5296 8676 5300 8732
rect 5236 8672 5300 8676
rect 10916 8732 10980 8736
rect 10916 8676 10920 8732
rect 10920 8676 10976 8732
rect 10976 8676 10980 8732
rect 10916 8672 10980 8676
rect 10996 8732 11060 8736
rect 10996 8676 11000 8732
rect 11000 8676 11056 8732
rect 11056 8676 11060 8732
rect 10996 8672 11060 8676
rect 11076 8732 11140 8736
rect 11076 8676 11080 8732
rect 11080 8676 11136 8732
rect 11136 8676 11140 8732
rect 11076 8672 11140 8676
rect 11156 8732 11220 8736
rect 11156 8676 11160 8732
rect 11160 8676 11216 8732
rect 11216 8676 11220 8732
rect 11156 8672 11220 8676
rect 11236 8732 11300 8736
rect 11236 8676 11240 8732
rect 11240 8676 11296 8732
rect 11296 8676 11300 8732
rect 11236 8672 11300 8676
rect 16916 8732 16980 8736
rect 16916 8676 16920 8732
rect 16920 8676 16976 8732
rect 16976 8676 16980 8732
rect 16916 8672 16980 8676
rect 16996 8732 17060 8736
rect 16996 8676 17000 8732
rect 17000 8676 17056 8732
rect 17056 8676 17060 8732
rect 16996 8672 17060 8676
rect 17076 8732 17140 8736
rect 17076 8676 17080 8732
rect 17080 8676 17136 8732
rect 17136 8676 17140 8732
rect 17076 8672 17140 8676
rect 17156 8732 17220 8736
rect 17156 8676 17160 8732
rect 17160 8676 17216 8732
rect 17216 8676 17220 8732
rect 17156 8672 17220 8676
rect 17236 8732 17300 8736
rect 17236 8676 17240 8732
rect 17240 8676 17296 8732
rect 17296 8676 17300 8732
rect 17236 8672 17300 8676
rect 22916 8732 22980 8736
rect 22916 8676 22920 8732
rect 22920 8676 22976 8732
rect 22976 8676 22980 8732
rect 22916 8672 22980 8676
rect 22996 8732 23060 8736
rect 22996 8676 23000 8732
rect 23000 8676 23056 8732
rect 23056 8676 23060 8732
rect 22996 8672 23060 8676
rect 23076 8732 23140 8736
rect 23076 8676 23080 8732
rect 23080 8676 23136 8732
rect 23136 8676 23140 8732
rect 23076 8672 23140 8676
rect 23156 8732 23220 8736
rect 23156 8676 23160 8732
rect 23160 8676 23216 8732
rect 23216 8676 23220 8732
rect 23156 8672 23220 8676
rect 23236 8732 23300 8736
rect 23236 8676 23240 8732
rect 23240 8676 23296 8732
rect 23296 8676 23300 8732
rect 23236 8672 23300 8676
rect 28916 8732 28980 8736
rect 28916 8676 28920 8732
rect 28920 8676 28976 8732
rect 28976 8676 28980 8732
rect 28916 8672 28980 8676
rect 28996 8732 29060 8736
rect 28996 8676 29000 8732
rect 29000 8676 29056 8732
rect 29056 8676 29060 8732
rect 28996 8672 29060 8676
rect 29076 8732 29140 8736
rect 29076 8676 29080 8732
rect 29080 8676 29136 8732
rect 29136 8676 29140 8732
rect 29076 8672 29140 8676
rect 29156 8732 29220 8736
rect 29156 8676 29160 8732
rect 29160 8676 29216 8732
rect 29216 8676 29220 8732
rect 29156 8672 29220 8676
rect 29236 8732 29300 8736
rect 29236 8676 29240 8732
rect 29240 8676 29296 8732
rect 29296 8676 29300 8732
rect 29236 8672 29300 8676
rect 4176 8188 4240 8192
rect 4176 8132 4180 8188
rect 4180 8132 4236 8188
rect 4236 8132 4240 8188
rect 4176 8128 4240 8132
rect 4256 8188 4320 8192
rect 4256 8132 4260 8188
rect 4260 8132 4316 8188
rect 4316 8132 4320 8188
rect 4256 8128 4320 8132
rect 4336 8188 4400 8192
rect 4336 8132 4340 8188
rect 4340 8132 4396 8188
rect 4396 8132 4400 8188
rect 4336 8128 4400 8132
rect 4416 8188 4480 8192
rect 4416 8132 4420 8188
rect 4420 8132 4476 8188
rect 4476 8132 4480 8188
rect 4416 8128 4480 8132
rect 4496 8188 4560 8192
rect 4496 8132 4500 8188
rect 4500 8132 4556 8188
rect 4556 8132 4560 8188
rect 4496 8128 4560 8132
rect 10176 8188 10240 8192
rect 10176 8132 10180 8188
rect 10180 8132 10236 8188
rect 10236 8132 10240 8188
rect 10176 8128 10240 8132
rect 10256 8188 10320 8192
rect 10256 8132 10260 8188
rect 10260 8132 10316 8188
rect 10316 8132 10320 8188
rect 10256 8128 10320 8132
rect 10336 8188 10400 8192
rect 10336 8132 10340 8188
rect 10340 8132 10396 8188
rect 10396 8132 10400 8188
rect 10336 8128 10400 8132
rect 10416 8188 10480 8192
rect 10416 8132 10420 8188
rect 10420 8132 10476 8188
rect 10476 8132 10480 8188
rect 10416 8128 10480 8132
rect 10496 8188 10560 8192
rect 10496 8132 10500 8188
rect 10500 8132 10556 8188
rect 10556 8132 10560 8188
rect 10496 8128 10560 8132
rect 16176 8188 16240 8192
rect 16176 8132 16180 8188
rect 16180 8132 16236 8188
rect 16236 8132 16240 8188
rect 16176 8128 16240 8132
rect 16256 8188 16320 8192
rect 16256 8132 16260 8188
rect 16260 8132 16316 8188
rect 16316 8132 16320 8188
rect 16256 8128 16320 8132
rect 16336 8188 16400 8192
rect 16336 8132 16340 8188
rect 16340 8132 16396 8188
rect 16396 8132 16400 8188
rect 16336 8128 16400 8132
rect 16416 8188 16480 8192
rect 16416 8132 16420 8188
rect 16420 8132 16476 8188
rect 16476 8132 16480 8188
rect 16416 8128 16480 8132
rect 16496 8188 16560 8192
rect 16496 8132 16500 8188
rect 16500 8132 16556 8188
rect 16556 8132 16560 8188
rect 16496 8128 16560 8132
rect 22176 8188 22240 8192
rect 22176 8132 22180 8188
rect 22180 8132 22236 8188
rect 22236 8132 22240 8188
rect 22176 8128 22240 8132
rect 22256 8188 22320 8192
rect 22256 8132 22260 8188
rect 22260 8132 22316 8188
rect 22316 8132 22320 8188
rect 22256 8128 22320 8132
rect 22336 8188 22400 8192
rect 22336 8132 22340 8188
rect 22340 8132 22396 8188
rect 22396 8132 22400 8188
rect 22336 8128 22400 8132
rect 22416 8188 22480 8192
rect 22416 8132 22420 8188
rect 22420 8132 22476 8188
rect 22476 8132 22480 8188
rect 22416 8128 22480 8132
rect 22496 8188 22560 8192
rect 22496 8132 22500 8188
rect 22500 8132 22556 8188
rect 22556 8132 22560 8188
rect 22496 8128 22560 8132
rect 28176 8188 28240 8192
rect 28176 8132 28180 8188
rect 28180 8132 28236 8188
rect 28236 8132 28240 8188
rect 28176 8128 28240 8132
rect 28256 8188 28320 8192
rect 28256 8132 28260 8188
rect 28260 8132 28316 8188
rect 28316 8132 28320 8188
rect 28256 8128 28320 8132
rect 28336 8188 28400 8192
rect 28336 8132 28340 8188
rect 28340 8132 28396 8188
rect 28396 8132 28400 8188
rect 28336 8128 28400 8132
rect 28416 8188 28480 8192
rect 28416 8132 28420 8188
rect 28420 8132 28476 8188
rect 28476 8132 28480 8188
rect 28416 8128 28480 8132
rect 28496 8188 28560 8192
rect 28496 8132 28500 8188
rect 28500 8132 28556 8188
rect 28556 8132 28560 8188
rect 28496 8128 28560 8132
rect 4916 7644 4980 7648
rect 4916 7588 4920 7644
rect 4920 7588 4976 7644
rect 4976 7588 4980 7644
rect 4916 7584 4980 7588
rect 4996 7644 5060 7648
rect 4996 7588 5000 7644
rect 5000 7588 5056 7644
rect 5056 7588 5060 7644
rect 4996 7584 5060 7588
rect 5076 7644 5140 7648
rect 5076 7588 5080 7644
rect 5080 7588 5136 7644
rect 5136 7588 5140 7644
rect 5076 7584 5140 7588
rect 5156 7644 5220 7648
rect 5156 7588 5160 7644
rect 5160 7588 5216 7644
rect 5216 7588 5220 7644
rect 5156 7584 5220 7588
rect 5236 7644 5300 7648
rect 5236 7588 5240 7644
rect 5240 7588 5296 7644
rect 5296 7588 5300 7644
rect 5236 7584 5300 7588
rect 10916 7644 10980 7648
rect 10916 7588 10920 7644
rect 10920 7588 10976 7644
rect 10976 7588 10980 7644
rect 10916 7584 10980 7588
rect 10996 7644 11060 7648
rect 10996 7588 11000 7644
rect 11000 7588 11056 7644
rect 11056 7588 11060 7644
rect 10996 7584 11060 7588
rect 11076 7644 11140 7648
rect 11076 7588 11080 7644
rect 11080 7588 11136 7644
rect 11136 7588 11140 7644
rect 11076 7584 11140 7588
rect 11156 7644 11220 7648
rect 11156 7588 11160 7644
rect 11160 7588 11216 7644
rect 11216 7588 11220 7644
rect 11156 7584 11220 7588
rect 11236 7644 11300 7648
rect 11236 7588 11240 7644
rect 11240 7588 11296 7644
rect 11296 7588 11300 7644
rect 11236 7584 11300 7588
rect 16916 7644 16980 7648
rect 16916 7588 16920 7644
rect 16920 7588 16976 7644
rect 16976 7588 16980 7644
rect 16916 7584 16980 7588
rect 16996 7644 17060 7648
rect 16996 7588 17000 7644
rect 17000 7588 17056 7644
rect 17056 7588 17060 7644
rect 16996 7584 17060 7588
rect 17076 7644 17140 7648
rect 17076 7588 17080 7644
rect 17080 7588 17136 7644
rect 17136 7588 17140 7644
rect 17076 7584 17140 7588
rect 17156 7644 17220 7648
rect 17156 7588 17160 7644
rect 17160 7588 17216 7644
rect 17216 7588 17220 7644
rect 17156 7584 17220 7588
rect 17236 7644 17300 7648
rect 17236 7588 17240 7644
rect 17240 7588 17296 7644
rect 17296 7588 17300 7644
rect 17236 7584 17300 7588
rect 22916 7644 22980 7648
rect 22916 7588 22920 7644
rect 22920 7588 22976 7644
rect 22976 7588 22980 7644
rect 22916 7584 22980 7588
rect 22996 7644 23060 7648
rect 22996 7588 23000 7644
rect 23000 7588 23056 7644
rect 23056 7588 23060 7644
rect 22996 7584 23060 7588
rect 23076 7644 23140 7648
rect 23076 7588 23080 7644
rect 23080 7588 23136 7644
rect 23136 7588 23140 7644
rect 23076 7584 23140 7588
rect 23156 7644 23220 7648
rect 23156 7588 23160 7644
rect 23160 7588 23216 7644
rect 23216 7588 23220 7644
rect 23156 7584 23220 7588
rect 23236 7644 23300 7648
rect 23236 7588 23240 7644
rect 23240 7588 23296 7644
rect 23296 7588 23300 7644
rect 23236 7584 23300 7588
rect 28916 7644 28980 7648
rect 28916 7588 28920 7644
rect 28920 7588 28976 7644
rect 28976 7588 28980 7644
rect 28916 7584 28980 7588
rect 28996 7644 29060 7648
rect 28996 7588 29000 7644
rect 29000 7588 29056 7644
rect 29056 7588 29060 7644
rect 28996 7584 29060 7588
rect 29076 7644 29140 7648
rect 29076 7588 29080 7644
rect 29080 7588 29136 7644
rect 29136 7588 29140 7644
rect 29076 7584 29140 7588
rect 29156 7644 29220 7648
rect 29156 7588 29160 7644
rect 29160 7588 29216 7644
rect 29216 7588 29220 7644
rect 29156 7584 29220 7588
rect 29236 7644 29300 7648
rect 29236 7588 29240 7644
rect 29240 7588 29296 7644
rect 29296 7588 29300 7644
rect 29236 7584 29300 7588
rect 4176 7100 4240 7104
rect 4176 7044 4180 7100
rect 4180 7044 4236 7100
rect 4236 7044 4240 7100
rect 4176 7040 4240 7044
rect 4256 7100 4320 7104
rect 4256 7044 4260 7100
rect 4260 7044 4316 7100
rect 4316 7044 4320 7100
rect 4256 7040 4320 7044
rect 4336 7100 4400 7104
rect 4336 7044 4340 7100
rect 4340 7044 4396 7100
rect 4396 7044 4400 7100
rect 4336 7040 4400 7044
rect 4416 7100 4480 7104
rect 4416 7044 4420 7100
rect 4420 7044 4476 7100
rect 4476 7044 4480 7100
rect 4416 7040 4480 7044
rect 4496 7100 4560 7104
rect 4496 7044 4500 7100
rect 4500 7044 4556 7100
rect 4556 7044 4560 7100
rect 4496 7040 4560 7044
rect 10176 7100 10240 7104
rect 10176 7044 10180 7100
rect 10180 7044 10236 7100
rect 10236 7044 10240 7100
rect 10176 7040 10240 7044
rect 10256 7100 10320 7104
rect 10256 7044 10260 7100
rect 10260 7044 10316 7100
rect 10316 7044 10320 7100
rect 10256 7040 10320 7044
rect 10336 7100 10400 7104
rect 10336 7044 10340 7100
rect 10340 7044 10396 7100
rect 10396 7044 10400 7100
rect 10336 7040 10400 7044
rect 10416 7100 10480 7104
rect 10416 7044 10420 7100
rect 10420 7044 10476 7100
rect 10476 7044 10480 7100
rect 10416 7040 10480 7044
rect 10496 7100 10560 7104
rect 10496 7044 10500 7100
rect 10500 7044 10556 7100
rect 10556 7044 10560 7100
rect 10496 7040 10560 7044
rect 16176 7100 16240 7104
rect 16176 7044 16180 7100
rect 16180 7044 16236 7100
rect 16236 7044 16240 7100
rect 16176 7040 16240 7044
rect 16256 7100 16320 7104
rect 16256 7044 16260 7100
rect 16260 7044 16316 7100
rect 16316 7044 16320 7100
rect 16256 7040 16320 7044
rect 16336 7100 16400 7104
rect 16336 7044 16340 7100
rect 16340 7044 16396 7100
rect 16396 7044 16400 7100
rect 16336 7040 16400 7044
rect 16416 7100 16480 7104
rect 16416 7044 16420 7100
rect 16420 7044 16476 7100
rect 16476 7044 16480 7100
rect 16416 7040 16480 7044
rect 16496 7100 16560 7104
rect 16496 7044 16500 7100
rect 16500 7044 16556 7100
rect 16556 7044 16560 7100
rect 16496 7040 16560 7044
rect 22176 7100 22240 7104
rect 22176 7044 22180 7100
rect 22180 7044 22236 7100
rect 22236 7044 22240 7100
rect 22176 7040 22240 7044
rect 22256 7100 22320 7104
rect 22256 7044 22260 7100
rect 22260 7044 22316 7100
rect 22316 7044 22320 7100
rect 22256 7040 22320 7044
rect 22336 7100 22400 7104
rect 22336 7044 22340 7100
rect 22340 7044 22396 7100
rect 22396 7044 22400 7100
rect 22336 7040 22400 7044
rect 22416 7100 22480 7104
rect 22416 7044 22420 7100
rect 22420 7044 22476 7100
rect 22476 7044 22480 7100
rect 22416 7040 22480 7044
rect 22496 7100 22560 7104
rect 22496 7044 22500 7100
rect 22500 7044 22556 7100
rect 22556 7044 22560 7100
rect 22496 7040 22560 7044
rect 28176 7100 28240 7104
rect 28176 7044 28180 7100
rect 28180 7044 28236 7100
rect 28236 7044 28240 7100
rect 28176 7040 28240 7044
rect 28256 7100 28320 7104
rect 28256 7044 28260 7100
rect 28260 7044 28316 7100
rect 28316 7044 28320 7100
rect 28256 7040 28320 7044
rect 28336 7100 28400 7104
rect 28336 7044 28340 7100
rect 28340 7044 28396 7100
rect 28396 7044 28400 7100
rect 28336 7040 28400 7044
rect 28416 7100 28480 7104
rect 28416 7044 28420 7100
rect 28420 7044 28476 7100
rect 28476 7044 28480 7100
rect 28416 7040 28480 7044
rect 28496 7100 28560 7104
rect 28496 7044 28500 7100
rect 28500 7044 28556 7100
rect 28556 7044 28560 7100
rect 28496 7040 28560 7044
rect 4916 6556 4980 6560
rect 4916 6500 4920 6556
rect 4920 6500 4976 6556
rect 4976 6500 4980 6556
rect 4916 6496 4980 6500
rect 4996 6556 5060 6560
rect 4996 6500 5000 6556
rect 5000 6500 5056 6556
rect 5056 6500 5060 6556
rect 4996 6496 5060 6500
rect 5076 6556 5140 6560
rect 5076 6500 5080 6556
rect 5080 6500 5136 6556
rect 5136 6500 5140 6556
rect 5076 6496 5140 6500
rect 5156 6556 5220 6560
rect 5156 6500 5160 6556
rect 5160 6500 5216 6556
rect 5216 6500 5220 6556
rect 5156 6496 5220 6500
rect 5236 6556 5300 6560
rect 5236 6500 5240 6556
rect 5240 6500 5296 6556
rect 5296 6500 5300 6556
rect 5236 6496 5300 6500
rect 10916 6556 10980 6560
rect 10916 6500 10920 6556
rect 10920 6500 10976 6556
rect 10976 6500 10980 6556
rect 10916 6496 10980 6500
rect 10996 6556 11060 6560
rect 10996 6500 11000 6556
rect 11000 6500 11056 6556
rect 11056 6500 11060 6556
rect 10996 6496 11060 6500
rect 11076 6556 11140 6560
rect 11076 6500 11080 6556
rect 11080 6500 11136 6556
rect 11136 6500 11140 6556
rect 11076 6496 11140 6500
rect 11156 6556 11220 6560
rect 11156 6500 11160 6556
rect 11160 6500 11216 6556
rect 11216 6500 11220 6556
rect 11156 6496 11220 6500
rect 11236 6556 11300 6560
rect 11236 6500 11240 6556
rect 11240 6500 11296 6556
rect 11296 6500 11300 6556
rect 11236 6496 11300 6500
rect 16916 6556 16980 6560
rect 16916 6500 16920 6556
rect 16920 6500 16976 6556
rect 16976 6500 16980 6556
rect 16916 6496 16980 6500
rect 16996 6556 17060 6560
rect 16996 6500 17000 6556
rect 17000 6500 17056 6556
rect 17056 6500 17060 6556
rect 16996 6496 17060 6500
rect 17076 6556 17140 6560
rect 17076 6500 17080 6556
rect 17080 6500 17136 6556
rect 17136 6500 17140 6556
rect 17076 6496 17140 6500
rect 17156 6556 17220 6560
rect 17156 6500 17160 6556
rect 17160 6500 17216 6556
rect 17216 6500 17220 6556
rect 17156 6496 17220 6500
rect 17236 6556 17300 6560
rect 17236 6500 17240 6556
rect 17240 6500 17296 6556
rect 17296 6500 17300 6556
rect 17236 6496 17300 6500
rect 22916 6556 22980 6560
rect 22916 6500 22920 6556
rect 22920 6500 22976 6556
rect 22976 6500 22980 6556
rect 22916 6496 22980 6500
rect 22996 6556 23060 6560
rect 22996 6500 23000 6556
rect 23000 6500 23056 6556
rect 23056 6500 23060 6556
rect 22996 6496 23060 6500
rect 23076 6556 23140 6560
rect 23076 6500 23080 6556
rect 23080 6500 23136 6556
rect 23136 6500 23140 6556
rect 23076 6496 23140 6500
rect 23156 6556 23220 6560
rect 23156 6500 23160 6556
rect 23160 6500 23216 6556
rect 23216 6500 23220 6556
rect 23156 6496 23220 6500
rect 23236 6556 23300 6560
rect 23236 6500 23240 6556
rect 23240 6500 23296 6556
rect 23296 6500 23300 6556
rect 23236 6496 23300 6500
rect 28916 6556 28980 6560
rect 28916 6500 28920 6556
rect 28920 6500 28976 6556
rect 28976 6500 28980 6556
rect 28916 6496 28980 6500
rect 28996 6556 29060 6560
rect 28996 6500 29000 6556
rect 29000 6500 29056 6556
rect 29056 6500 29060 6556
rect 28996 6496 29060 6500
rect 29076 6556 29140 6560
rect 29076 6500 29080 6556
rect 29080 6500 29136 6556
rect 29136 6500 29140 6556
rect 29076 6496 29140 6500
rect 29156 6556 29220 6560
rect 29156 6500 29160 6556
rect 29160 6500 29216 6556
rect 29216 6500 29220 6556
rect 29156 6496 29220 6500
rect 29236 6556 29300 6560
rect 29236 6500 29240 6556
rect 29240 6500 29296 6556
rect 29296 6500 29300 6556
rect 29236 6496 29300 6500
rect 4176 6012 4240 6016
rect 4176 5956 4180 6012
rect 4180 5956 4236 6012
rect 4236 5956 4240 6012
rect 4176 5952 4240 5956
rect 4256 6012 4320 6016
rect 4256 5956 4260 6012
rect 4260 5956 4316 6012
rect 4316 5956 4320 6012
rect 4256 5952 4320 5956
rect 4336 6012 4400 6016
rect 4336 5956 4340 6012
rect 4340 5956 4396 6012
rect 4396 5956 4400 6012
rect 4336 5952 4400 5956
rect 4416 6012 4480 6016
rect 4416 5956 4420 6012
rect 4420 5956 4476 6012
rect 4476 5956 4480 6012
rect 4416 5952 4480 5956
rect 4496 6012 4560 6016
rect 4496 5956 4500 6012
rect 4500 5956 4556 6012
rect 4556 5956 4560 6012
rect 4496 5952 4560 5956
rect 10176 6012 10240 6016
rect 10176 5956 10180 6012
rect 10180 5956 10236 6012
rect 10236 5956 10240 6012
rect 10176 5952 10240 5956
rect 10256 6012 10320 6016
rect 10256 5956 10260 6012
rect 10260 5956 10316 6012
rect 10316 5956 10320 6012
rect 10256 5952 10320 5956
rect 10336 6012 10400 6016
rect 10336 5956 10340 6012
rect 10340 5956 10396 6012
rect 10396 5956 10400 6012
rect 10336 5952 10400 5956
rect 10416 6012 10480 6016
rect 10416 5956 10420 6012
rect 10420 5956 10476 6012
rect 10476 5956 10480 6012
rect 10416 5952 10480 5956
rect 10496 6012 10560 6016
rect 10496 5956 10500 6012
rect 10500 5956 10556 6012
rect 10556 5956 10560 6012
rect 10496 5952 10560 5956
rect 16176 6012 16240 6016
rect 16176 5956 16180 6012
rect 16180 5956 16236 6012
rect 16236 5956 16240 6012
rect 16176 5952 16240 5956
rect 16256 6012 16320 6016
rect 16256 5956 16260 6012
rect 16260 5956 16316 6012
rect 16316 5956 16320 6012
rect 16256 5952 16320 5956
rect 16336 6012 16400 6016
rect 16336 5956 16340 6012
rect 16340 5956 16396 6012
rect 16396 5956 16400 6012
rect 16336 5952 16400 5956
rect 16416 6012 16480 6016
rect 16416 5956 16420 6012
rect 16420 5956 16476 6012
rect 16476 5956 16480 6012
rect 16416 5952 16480 5956
rect 16496 6012 16560 6016
rect 16496 5956 16500 6012
rect 16500 5956 16556 6012
rect 16556 5956 16560 6012
rect 16496 5952 16560 5956
rect 22176 6012 22240 6016
rect 22176 5956 22180 6012
rect 22180 5956 22236 6012
rect 22236 5956 22240 6012
rect 22176 5952 22240 5956
rect 22256 6012 22320 6016
rect 22256 5956 22260 6012
rect 22260 5956 22316 6012
rect 22316 5956 22320 6012
rect 22256 5952 22320 5956
rect 22336 6012 22400 6016
rect 22336 5956 22340 6012
rect 22340 5956 22396 6012
rect 22396 5956 22400 6012
rect 22336 5952 22400 5956
rect 22416 6012 22480 6016
rect 22416 5956 22420 6012
rect 22420 5956 22476 6012
rect 22476 5956 22480 6012
rect 22416 5952 22480 5956
rect 22496 6012 22560 6016
rect 22496 5956 22500 6012
rect 22500 5956 22556 6012
rect 22556 5956 22560 6012
rect 22496 5952 22560 5956
rect 28176 6012 28240 6016
rect 28176 5956 28180 6012
rect 28180 5956 28236 6012
rect 28236 5956 28240 6012
rect 28176 5952 28240 5956
rect 28256 6012 28320 6016
rect 28256 5956 28260 6012
rect 28260 5956 28316 6012
rect 28316 5956 28320 6012
rect 28256 5952 28320 5956
rect 28336 6012 28400 6016
rect 28336 5956 28340 6012
rect 28340 5956 28396 6012
rect 28396 5956 28400 6012
rect 28336 5952 28400 5956
rect 28416 6012 28480 6016
rect 28416 5956 28420 6012
rect 28420 5956 28476 6012
rect 28476 5956 28480 6012
rect 28416 5952 28480 5956
rect 28496 6012 28560 6016
rect 28496 5956 28500 6012
rect 28500 5956 28556 6012
rect 28556 5956 28560 6012
rect 28496 5952 28560 5956
rect 4916 5468 4980 5472
rect 4916 5412 4920 5468
rect 4920 5412 4976 5468
rect 4976 5412 4980 5468
rect 4916 5408 4980 5412
rect 4996 5468 5060 5472
rect 4996 5412 5000 5468
rect 5000 5412 5056 5468
rect 5056 5412 5060 5468
rect 4996 5408 5060 5412
rect 5076 5468 5140 5472
rect 5076 5412 5080 5468
rect 5080 5412 5136 5468
rect 5136 5412 5140 5468
rect 5076 5408 5140 5412
rect 5156 5468 5220 5472
rect 5156 5412 5160 5468
rect 5160 5412 5216 5468
rect 5216 5412 5220 5468
rect 5156 5408 5220 5412
rect 5236 5468 5300 5472
rect 5236 5412 5240 5468
rect 5240 5412 5296 5468
rect 5296 5412 5300 5468
rect 5236 5408 5300 5412
rect 10916 5468 10980 5472
rect 10916 5412 10920 5468
rect 10920 5412 10976 5468
rect 10976 5412 10980 5468
rect 10916 5408 10980 5412
rect 10996 5468 11060 5472
rect 10996 5412 11000 5468
rect 11000 5412 11056 5468
rect 11056 5412 11060 5468
rect 10996 5408 11060 5412
rect 11076 5468 11140 5472
rect 11076 5412 11080 5468
rect 11080 5412 11136 5468
rect 11136 5412 11140 5468
rect 11076 5408 11140 5412
rect 11156 5468 11220 5472
rect 11156 5412 11160 5468
rect 11160 5412 11216 5468
rect 11216 5412 11220 5468
rect 11156 5408 11220 5412
rect 11236 5468 11300 5472
rect 11236 5412 11240 5468
rect 11240 5412 11296 5468
rect 11296 5412 11300 5468
rect 11236 5408 11300 5412
rect 16916 5468 16980 5472
rect 16916 5412 16920 5468
rect 16920 5412 16976 5468
rect 16976 5412 16980 5468
rect 16916 5408 16980 5412
rect 16996 5468 17060 5472
rect 16996 5412 17000 5468
rect 17000 5412 17056 5468
rect 17056 5412 17060 5468
rect 16996 5408 17060 5412
rect 17076 5468 17140 5472
rect 17076 5412 17080 5468
rect 17080 5412 17136 5468
rect 17136 5412 17140 5468
rect 17076 5408 17140 5412
rect 17156 5468 17220 5472
rect 17156 5412 17160 5468
rect 17160 5412 17216 5468
rect 17216 5412 17220 5468
rect 17156 5408 17220 5412
rect 17236 5468 17300 5472
rect 17236 5412 17240 5468
rect 17240 5412 17296 5468
rect 17296 5412 17300 5468
rect 17236 5408 17300 5412
rect 22916 5468 22980 5472
rect 22916 5412 22920 5468
rect 22920 5412 22976 5468
rect 22976 5412 22980 5468
rect 22916 5408 22980 5412
rect 22996 5468 23060 5472
rect 22996 5412 23000 5468
rect 23000 5412 23056 5468
rect 23056 5412 23060 5468
rect 22996 5408 23060 5412
rect 23076 5468 23140 5472
rect 23076 5412 23080 5468
rect 23080 5412 23136 5468
rect 23136 5412 23140 5468
rect 23076 5408 23140 5412
rect 23156 5468 23220 5472
rect 23156 5412 23160 5468
rect 23160 5412 23216 5468
rect 23216 5412 23220 5468
rect 23156 5408 23220 5412
rect 23236 5468 23300 5472
rect 23236 5412 23240 5468
rect 23240 5412 23296 5468
rect 23296 5412 23300 5468
rect 23236 5408 23300 5412
rect 28916 5468 28980 5472
rect 28916 5412 28920 5468
rect 28920 5412 28976 5468
rect 28976 5412 28980 5468
rect 28916 5408 28980 5412
rect 28996 5468 29060 5472
rect 28996 5412 29000 5468
rect 29000 5412 29056 5468
rect 29056 5412 29060 5468
rect 28996 5408 29060 5412
rect 29076 5468 29140 5472
rect 29076 5412 29080 5468
rect 29080 5412 29136 5468
rect 29136 5412 29140 5468
rect 29076 5408 29140 5412
rect 29156 5468 29220 5472
rect 29156 5412 29160 5468
rect 29160 5412 29216 5468
rect 29216 5412 29220 5468
rect 29156 5408 29220 5412
rect 29236 5468 29300 5472
rect 29236 5412 29240 5468
rect 29240 5412 29296 5468
rect 29296 5412 29300 5468
rect 29236 5408 29300 5412
rect 4176 4924 4240 4928
rect 4176 4868 4180 4924
rect 4180 4868 4236 4924
rect 4236 4868 4240 4924
rect 4176 4864 4240 4868
rect 4256 4924 4320 4928
rect 4256 4868 4260 4924
rect 4260 4868 4316 4924
rect 4316 4868 4320 4924
rect 4256 4864 4320 4868
rect 4336 4924 4400 4928
rect 4336 4868 4340 4924
rect 4340 4868 4396 4924
rect 4396 4868 4400 4924
rect 4336 4864 4400 4868
rect 4416 4924 4480 4928
rect 4416 4868 4420 4924
rect 4420 4868 4476 4924
rect 4476 4868 4480 4924
rect 4416 4864 4480 4868
rect 4496 4924 4560 4928
rect 4496 4868 4500 4924
rect 4500 4868 4556 4924
rect 4556 4868 4560 4924
rect 4496 4864 4560 4868
rect 10176 4924 10240 4928
rect 10176 4868 10180 4924
rect 10180 4868 10236 4924
rect 10236 4868 10240 4924
rect 10176 4864 10240 4868
rect 10256 4924 10320 4928
rect 10256 4868 10260 4924
rect 10260 4868 10316 4924
rect 10316 4868 10320 4924
rect 10256 4864 10320 4868
rect 10336 4924 10400 4928
rect 10336 4868 10340 4924
rect 10340 4868 10396 4924
rect 10396 4868 10400 4924
rect 10336 4864 10400 4868
rect 10416 4924 10480 4928
rect 10416 4868 10420 4924
rect 10420 4868 10476 4924
rect 10476 4868 10480 4924
rect 10416 4864 10480 4868
rect 10496 4924 10560 4928
rect 10496 4868 10500 4924
rect 10500 4868 10556 4924
rect 10556 4868 10560 4924
rect 10496 4864 10560 4868
rect 16176 4924 16240 4928
rect 16176 4868 16180 4924
rect 16180 4868 16236 4924
rect 16236 4868 16240 4924
rect 16176 4864 16240 4868
rect 16256 4924 16320 4928
rect 16256 4868 16260 4924
rect 16260 4868 16316 4924
rect 16316 4868 16320 4924
rect 16256 4864 16320 4868
rect 16336 4924 16400 4928
rect 16336 4868 16340 4924
rect 16340 4868 16396 4924
rect 16396 4868 16400 4924
rect 16336 4864 16400 4868
rect 16416 4924 16480 4928
rect 16416 4868 16420 4924
rect 16420 4868 16476 4924
rect 16476 4868 16480 4924
rect 16416 4864 16480 4868
rect 16496 4924 16560 4928
rect 16496 4868 16500 4924
rect 16500 4868 16556 4924
rect 16556 4868 16560 4924
rect 16496 4864 16560 4868
rect 22176 4924 22240 4928
rect 22176 4868 22180 4924
rect 22180 4868 22236 4924
rect 22236 4868 22240 4924
rect 22176 4864 22240 4868
rect 22256 4924 22320 4928
rect 22256 4868 22260 4924
rect 22260 4868 22316 4924
rect 22316 4868 22320 4924
rect 22256 4864 22320 4868
rect 22336 4924 22400 4928
rect 22336 4868 22340 4924
rect 22340 4868 22396 4924
rect 22396 4868 22400 4924
rect 22336 4864 22400 4868
rect 22416 4924 22480 4928
rect 22416 4868 22420 4924
rect 22420 4868 22476 4924
rect 22476 4868 22480 4924
rect 22416 4864 22480 4868
rect 22496 4924 22560 4928
rect 22496 4868 22500 4924
rect 22500 4868 22556 4924
rect 22556 4868 22560 4924
rect 22496 4864 22560 4868
rect 28176 4924 28240 4928
rect 28176 4868 28180 4924
rect 28180 4868 28236 4924
rect 28236 4868 28240 4924
rect 28176 4864 28240 4868
rect 28256 4924 28320 4928
rect 28256 4868 28260 4924
rect 28260 4868 28316 4924
rect 28316 4868 28320 4924
rect 28256 4864 28320 4868
rect 28336 4924 28400 4928
rect 28336 4868 28340 4924
rect 28340 4868 28396 4924
rect 28396 4868 28400 4924
rect 28336 4864 28400 4868
rect 28416 4924 28480 4928
rect 28416 4868 28420 4924
rect 28420 4868 28476 4924
rect 28476 4868 28480 4924
rect 28416 4864 28480 4868
rect 28496 4924 28560 4928
rect 28496 4868 28500 4924
rect 28500 4868 28556 4924
rect 28556 4868 28560 4924
rect 28496 4864 28560 4868
rect 4916 4380 4980 4384
rect 4916 4324 4920 4380
rect 4920 4324 4976 4380
rect 4976 4324 4980 4380
rect 4916 4320 4980 4324
rect 4996 4380 5060 4384
rect 4996 4324 5000 4380
rect 5000 4324 5056 4380
rect 5056 4324 5060 4380
rect 4996 4320 5060 4324
rect 5076 4380 5140 4384
rect 5076 4324 5080 4380
rect 5080 4324 5136 4380
rect 5136 4324 5140 4380
rect 5076 4320 5140 4324
rect 5156 4380 5220 4384
rect 5156 4324 5160 4380
rect 5160 4324 5216 4380
rect 5216 4324 5220 4380
rect 5156 4320 5220 4324
rect 5236 4380 5300 4384
rect 5236 4324 5240 4380
rect 5240 4324 5296 4380
rect 5296 4324 5300 4380
rect 5236 4320 5300 4324
rect 10916 4380 10980 4384
rect 10916 4324 10920 4380
rect 10920 4324 10976 4380
rect 10976 4324 10980 4380
rect 10916 4320 10980 4324
rect 10996 4380 11060 4384
rect 10996 4324 11000 4380
rect 11000 4324 11056 4380
rect 11056 4324 11060 4380
rect 10996 4320 11060 4324
rect 11076 4380 11140 4384
rect 11076 4324 11080 4380
rect 11080 4324 11136 4380
rect 11136 4324 11140 4380
rect 11076 4320 11140 4324
rect 11156 4380 11220 4384
rect 11156 4324 11160 4380
rect 11160 4324 11216 4380
rect 11216 4324 11220 4380
rect 11156 4320 11220 4324
rect 11236 4380 11300 4384
rect 11236 4324 11240 4380
rect 11240 4324 11296 4380
rect 11296 4324 11300 4380
rect 11236 4320 11300 4324
rect 16916 4380 16980 4384
rect 16916 4324 16920 4380
rect 16920 4324 16976 4380
rect 16976 4324 16980 4380
rect 16916 4320 16980 4324
rect 16996 4380 17060 4384
rect 16996 4324 17000 4380
rect 17000 4324 17056 4380
rect 17056 4324 17060 4380
rect 16996 4320 17060 4324
rect 17076 4380 17140 4384
rect 17076 4324 17080 4380
rect 17080 4324 17136 4380
rect 17136 4324 17140 4380
rect 17076 4320 17140 4324
rect 17156 4380 17220 4384
rect 17156 4324 17160 4380
rect 17160 4324 17216 4380
rect 17216 4324 17220 4380
rect 17156 4320 17220 4324
rect 17236 4380 17300 4384
rect 17236 4324 17240 4380
rect 17240 4324 17296 4380
rect 17296 4324 17300 4380
rect 17236 4320 17300 4324
rect 22916 4380 22980 4384
rect 22916 4324 22920 4380
rect 22920 4324 22976 4380
rect 22976 4324 22980 4380
rect 22916 4320 22980 4324
rect 22996 4380 23060 4384
rect 22996 4324 23000 4380
rect 23000 4324 23056 4380
rect 23056 4324 23060 4380
rect 22996 4320 23060 4324
rect 23076 4380 23140 4384
rect 23076 4324 23080 4380
rect 23080 4324 23136 4380
rect 23136 4324 23140 4380
rect 23076 4320 23140 4324
rect 23156 4380 23220 4384
rect 23156 4324 23160 4380
rect 23160 4324 23216 4380
rect 23216 4324 23220 4380
rect 23156 4320 23220 4324
rect 23236 4380 23300 4384
rect 23236 4324 23240 4380
rect 23240 4324 23296 4380
rect 23296 4324 23300 4380
rect 23236 4320 23300 4324
rect 28916 4380 28980 4384
rect 28916 4324 28920 4380
rect 28920 4324 28976 4380
rect 28976 4324 28980 4380
rect 28916 4320 28980 4324
rect 28996 4380 29060 4384
rect 28996 4324 29000 4380
rect 29000 4324 29056 4380
rect 29056 4324 29060 4380
rect 28996 4320 29060 4324
rect 29076 4380 29140 4384
rect 29076 4324 29080 4380
rect 29080 4324 29136 4380
rect 29136 4324 29140 4380
rect 29076 4320 29140 4324
rect 29156 4380 29220 4384
rect 29156 4324 29160 4380
rect 29160 4324 29216 4380
rect 29216 4324 29220 4380
rect 29156 4320 29220 4324
rect 29236 4380 29300 4384
rect 29236 4324 29240 4380
rect 29240 4324 29296 4380
rect 29296 4324 29300 4380
rect 29236 4320 29300 4324
rect 4176 3836 4240 3840
rect 4176 3780 4180 3836
rect 4180 3780 4236 3836
rect 4236 3780 4240 3836
rect 4176 3776 4240 3780
rect 4256 3836 4320 3840
rect 4256 3780 4260 3836
rect 4260 3780 4316 3836
rect 4316 3780 4320 3836
rect 4256 3776 4320 3780
rect 4336 3836 4400 3840
rect 4336 3780 4340 3836
rect 4340 3780 4396 3836
rect 4396 3780 4400 3836
rect 4336 3776 4400 3780
rect 4416 3836 4480 3840
rect 4416 3780 4420 3836
rect 4420 3780 4476 3836
rect 4476 3780 4480 3836
rect 4416 3776 4480 3780
rect 4496 3836 4560 3840
rect 4496 3780 4500 3836
rect 4500 3780 4556 3836
rect 4556 3780 4560 3836
rect 4496 3776 4560 3780
rect 10176 3836 10240 3840
rect 10176 3780 10180 3836
rect 10180 3780 10236 3836
rect 10236 3780 10240 3836
rect 10176 3776 10240 3780
rect 10256 3836 10320 3840
rect 10256 3780 10260 3836
rect 10260 3780 10316 3836
rect 10316 3780 10320 3836
rect 10256 3776 10320 3780
rect 10336 3836 10400 3840
rect 10336 3780 10340 3836
rect 10340 3780 10396 3836
rect 10396 3780 10400 3836
rect 10336 3776 10400 3780
rect 10416 3836 10480 3840
rect 10416 3780 10420 3836
rect 10420 3780 10476 3836
rect 10476 3780 10480 3836
rect 10416 3776 10480 3780
rect 10496 3836 10560 3840
rect 10496 3780 10500 3836
rect 10500 3780 10556 3836
rect 10556 3780 10560 3836
rect 10496 3776 10560 3780
rect 16176 3836 16240 3840
rect 16176 3780 16180 3836
rect 16180 3780 16236 3836
rect 16236 3780 16240 3836
rect 16176 3776 16240 3780
rect 16256 3836 16320 3840
rect 16256 3780 16260 3836
rect 16260 3780 16316 3836
rect 16316 3780 16320 3836
rect 16256 3776 16320 3780
rect 16336 3836 16400 3840
rect 16336 3780 16340 3836
rect 16340 3780 16396 3836
rect 16396 3780 16400 3836
rect 16336 3776 16400 3780
rect 16416 3836 16480 3840
rect 16416 3780 16420 3836
rect 16420 3780 16476 3836
rect 16476 3780 16480 3836
rect 16416 3776 16480 3780
rect 16496 3836 16560 3840
rect 16496 3780 16500 3836
rect 16500 3780 16556 3836
rect 16556 3780 16560 3836
rect 16496 3776 16560 3780
rect 22176 3836 22240 3840
rect 22176 3780 22180 3836
rect 22180 3780 22236 3836
rect 22236 3780 22240 3836
rect 22176 3776 22240 3780
rect 22256 3836 22320 3840
rect 22256 3780 22260 3836
rect 22260 3780 22316 3836
rect 22316 3780 22320 3836
rect 22256 3776 22320 3780
rect 22336 3836 22400 3840
rect 22336 3780 22340 3836
rect 22340 3780 22396 3836
rect 22396 3780 22400 3836
rect 22336 3776 22400 3780
rect 22416 3836 22480 3840
rect 22416 3780 22420 3836
rect 22420 3780 22476 3836
rect 22476 3780 22480 3836
rect 22416 3776 22480 3780
rect 22496 3836 22560 3840
rect 22496 3780 22500 3836
rect 22500 3780 22556 3836
rect 22556 3780 22560 3836
rect 22496 3776 22560 3780
rect 28176 3836 28240 3840
rect 28176 3780 28180 3836
rect 28180 3780 28236 3836
rect 28236 3780 28240 3836
rect 28176 3776 28240 3780
rect 28256 3836 28320 3840
rect 28256 3780 28260 3836
rect 28260 3780 28316 3836
rect 28316 3780 28320 3836
rect 28256 3776 28320 3780
rect 28336 3836 28400 3840
rect 28336 3780 28340 3836
rect 28340 3780 28396 3836
rect 28396 3780 28400 3836
rect 28336 3776 28400 3780
rect 28416 3836 28480 3840
rect 28416 3780 28420 3836
rect 28420 3780 28476 3836
rect 28476 3780 28480 3836
rect 28416 3776 28480 3780
rect 28496 3836 28560 3840
rect 28496 3780 28500 3836
rect 28500 3780 28556 3836
rect 28556 3780 28560 3836
rect 28496 3776 28560 3780
rect 4916 3292 4980 3296
rect 4916 3236 4920 3292
rect 4920 3236 4976 3292
rect 4976 3236 4980 3292
rect 4916 3232 4980 3236
rect 4996 3292 5060 3296
rect 4996 3236 5000 3292
rect 5000 3236 5056 3292
rect 5056 3236 5060 3292
rect 4996 3232 5060 3236
rect 5076 3292 5140 3296
rect 5076 3236 5080 3292
rect 5080 3236 5136 3292
rect 5136 3236 5140 3292
rect 5076 3232 5140 3236
rect 5156 3292 5220 3296
rect 5156 3236 5160 3292
rect 5160 3236 5216 3292
rect 5216 3236 5220 3292
rect 5156 3232 5220 3236
rect 5236 3292 5300 3296
rect 5236 3236 5240 3292
rect 5240 3236 5296 3292
rect 5296 3236 5300 3292
rect 5236 3232 5300 3236
rect 10916 3292 10980 3296
rect 10916 3236 10920 3292
rect 10920 3236 10976 3292
rect 10976 3236 10980 3292
rect 10916 3232 10980 3236
rect 10996 3292 11060 3296
rect 10996 3236 11000 3292
rect 11000 3236 11056 3292
rect 11056 3236 11060 3292
rect 10996 3232 11060 3236
rect 11076 3292 11140 3296
rect 11076 3236 11080 3292
rect 11080 3236 11136 3292
rect 11136 3236 11140 3292
rect 11076 3232 11140 3236
rect 11156 3292 11220 3296
rect 11156 3236 11160 3292
rect 11160 3236 11216 3292
rect 11216 3236 11220 3292
rect 11156 3232 11220 3236
rect 11236 3292 11300 3296
rect 11236 3236 11240 3292
rect 11240 3236 11296 3292
rect 11296 3236 11300 3292
rect 11236 3232 11300 3236
rect 16916 3292 16980 3296
rect 16916 3236 16920 3292
rect 16920 3236 16976 3292
rect 16976 3236 16980 3292
rect 16916 3232 16980 3236
rect 16996 3292 17060 3296
rect 16996 3236 17000 3292
rect 17000 3236 17056 3292
rect 17056 3236 17060 3292
rect 16996 3232 17060 3236
rect 17076 3292 17140 3296
rect 17076 3236 17080 3292
rect 17080 3236 17136 3292
rect 17136 3236 17140 3292
rect 17076 3232 17140 3236
rect 17156 3292 17220 3296
rect 17156 3236 17160 3292
rect 17160 3236 17216 3292
rect 17216 3236 17220 3292
rect 17156 3232 17220 3236
rect 17236 3292 17300 3296
rect 17236 3236 17240 3292
rect 17240 3236 17296 3292
rect 17296 3236 17300 3292
rect 17236 3232 17300 3236
rect 22916 3292 22980 3296
rect 22916 3236 22920 3292
rect 22920 3236 22976 3292
rect 22976 3236 22980 3292
rect 22916 3232 22980 3236
rect 22996 3292 23060 3296
rect 22996 3236 23000 3292
rect 23000 3236 23056 3292
rect 23056 3236 23060 3292
rect 22996 3232 23060 3236
rect 23076 3292 23140 3296
rect 23076 3236 23080 3292
rect 23080 3236 23136 3292
rect 23136 3236 23140 3292
rect 23076 3232 23140 3236
rect 23156 3292 23220 3296
rect 23156 3236 23160 3292
rect 23160 3236 23216 3292
rect 23216 3236 23220 3292
rect 23156 3232 23220 3236
rect 23236 3292 23300 3296
rect 23236 3236 23240 3292
rect 23240 3236 23296 3292
rect 23296 3236 23300 3292
rect 23236 3232 23300 3236
rect 28916 3292 28980 3296
rect 28916 3236 28920 3292
rect 28920 3236 28976 3292
rect 28976 3236 28980 3292
rect 28916 3232 28980 3236
rect 28996 3292 29060 3296
rect 28996 3236 29000 3292
rect 29000 3236 29056 3292
rect 29056 3236 29060 3292
rect 28996 3232 29060 3236
rect 29076 3292 29140 3296
rect 29076 3236 29080 3292
rect 29080 3236 29136 3292
rect 29136 3236 29140 3292
rect 29076 3232 29140 3236
rect 29156 3292 29220 3296
rect 29156 3236 29160 3292
rect 29160 3236 29216 3292
rect 29216 3236 29220 3292
rect 29156 3232 29220 3236
rect 29236 3292 29300 3296
rect 29236 3236 29240 3292
rect 29240 3236 29296 3292
rect 29296 3236 29300 3292
rect 29236 3232 29300 3236
rect 4176 2748 4240 2752
rect 4176 2692 4180 2748
rect 4180 2692 4236 2748
rect 4236 2692 4240 2748
rect 4176 2688 4240 2692
rect 4256 2748 4320 2752
rect 4256 2692 4260 2748
rect 4260 2692 4316 2748
rect 4316 2692 4320 2748
rect 4256 2688 4320 2692
rect 4336 2748 4400 2752
rect 4336 2692 4340 2748
rect 4340 2692 4396 2748
rect 4396 2692 4400 2748
rect 4336 2688 4400 2692
rect 4416 2748 4480 2752
rect 4416 2692 4420 2748
rect 4420 2692 4476 2748
rect 4476 2692 4480 2748
rect 4416 2688 4480 2692
rect 4496 2748 4560 2752
rect 4496 2692 4500 2748
rect 4500 2692 4556 2748
rect 4556 2692 4560 2748
rect 4496 2688 4560 2692
rect 10176 2748 10240 2752
rect 10176 2692 10180 2748
rect 10180 2692 10236 2748
rect 10236 2692 10240 2748
rect 10176 2688 10240 2692
rect 10256 2748 10320 2752
rect 10256 2692 10260 2748
rect 10260 2692 10316 2748
rect 10316 2692 10320 2748
rect 10256 2688 10320 2692
rect 10336 2748 10400 2752
rect 10336 2692 10340 2748
rect 10340 2692 10396 2748
rect 10396 2692 10400 2748
rect 10336 2688 10400 2692
rect 10416 2748 10480 2752
rect 10416 2692 10420 2748
rect 10420 2692 10476 2748
rect 10476 2692 10480 2748
rect 10416 2688 10480 2692
rect 10496 2748 10560 2752
rect 10496 2692 10500 2748
rect 10500 2692 10556 2748
rect 10556 2692 10560 2748
rect 10496 2688 10560 2692
rect 16176 2748 16240 2752
rect 16176 2692 16180 2748
rect 16180 2692 16236 2748
rect 16236 2692 16240 2748
rect 16176 2688 16240 2692
rect 16256 2748 16320 2752
rect 16256 2692 16260 2748
rect 16260 2692 16316 2748
rect 16316 2692 16320 2748
rect 16256 2688 16320 2692
rect 16336 2748 16400 2752
rect 16336 2692 16340 2748
rect 16340 2692 16396 2748
rect 16396 2692 16400 2748
rect 16336 2688 16400 2692
rect 16416 2748 16480 2752
rect 16416 2692 16420 2748
rect 16420 2692 16476 2748
rect 16476 2692 16480 2748
rect 16416 2688 16480 2692
rect 16496 2748 16560 2752
rect 16496 2692 16500 2748
rect 16500 2692 16556 2748
rect 16556 2692 16560 2748
rect 16496 2688 16560 2692
rect 22176 2748 22240 2752
rect 22176 2692 22180 2748
rect 22180 2692 22236 2748
rect 22236 2692 22240 2748
rect 22176 2688 22240 2692
rect 22256 2748 22320 2752
rect 22256 2692 22260 2748
rect 22260 2692 22316 2748
rect 22316 2692 22320 2748
rect 22256 2688 22320 2692
rect 22336 2748 22400 2752
rect 22336 2692 22340 2748
rect 22340 2692 22396 2748
rect 22396 2692 22400 2748
rect 22336 2688 22400 2692
rect 22416 2748 22480 2752
rect 22416 2692 22420 2748
rect 22420 2692 22476 2748
rect 22476 2692 22480 2748
rect 22416 2688 22480 2692
rect 22496 2748 22560 2752
rect 22496 2692 22500 2748
rect 22500 2692 22556 2748
rect 22556 2692 22560 2748
rect 22496 2688 22560 2692
rect 28176 2748 28240 2752
rect 28176 2692 28180 2748
rect 28180 2692 28236 2748
rect 28236 2692 28240 2748
rect 28176 2688 28240 2692
rect 28256 2748 28320 2752
rect 28256 2692 28260 2748
rect 28260 2692 28316 2748
rect 28316 2692 28320 2748
rect 28256 2688 28320 2692
rect 28336 2748 28400 2752
rect 28336 2692 28340 2748
rect 28340 2692 28396 2748
rect 28396 2692 28400 2748
rect 28336 2688 28400 2692
rect 28416 2748 28480 2752
rect 28416 2692 28420 2748
rect 28420 2692 28476 2748
rect 28476 2692 28480 2748
rect 28416 2688 28480 2692
rect 28496 2748 28560 2752
rect 28496 2692 28500 2748
rect 28500 2692 28556 2748
rect 28556 2692 28560 2748
rect 28496 2688 28560 2692
rect 4916 2204 4980 2208
rect 4916 2148 4920 2204
rect 4920 2148 4976 2204
rect 4976 2148 4980 2204
rect 4916 2144 4980 2148
rect 4996 2204 5060 2208
rect 4996 2148 5000 2204
rect 5000 2148 5056 2204
rect 5056 2148 5060 2204
rect 4996 2144 5060 2148
rect 5076 2204 5140 2208
rect 5076 2148 5080 2204
rect 5080 2148 5136 2204
rect 5136 2148 5140 2204
rect 5076 2144 5140 2148
rect 5156 2204 5220 2208
rect 5156 2148 5160 2204
rect 5160 2148 5216 2204
rect 5216 2148 5220 2204
rect 5156 2144 5220 2148
rect 5236 2204 5300 2208
rect 5236 2148 5240 2204
rect 5240 2148 5296 2204
rect 5296 2148 5300 2204
rect 5236 2144 5300 2148
rect 10916 2204 10980 2208
rect 10916 2148 10920 2204
rect 10920 2148 10976 2204
rect 10976 2148 10980 2204
rect 10916 2144 10980 2148
rect 10996 2204 11060 2208
rect 10996 2148 11000 2204
rect 11000 2148 11056 2204
rect 11056 2148 11060 2204
rect 10996 2144 11060 2148
rect 11076 2204 11140 2208
rect 11076 2148 11080 2204
rect 11080 2148 11136 2204
rect 11136 2148 11140 2204
rect 11076 2144 11140 2148
rect 11156 2204 11220 2208
rect 11156 2148 11160 2204
rect 11160 2148 11216 2204
rect 11216 2148 11220 2204
rect 11156 2144 11220 2148
rect 11236 2204 11300 2208
rect 11236 2148 11240 2204
rect 11240 2148 11296 2204
rect 11296 2148 11300 2204
rect 11236 2144 11300 2148
rect 16916 2204 16980 2208
rect 16916 2148 16920 2204
rect 16920 2148 16976 2204
rect 16976 2148 16980 2204
rect 16916 2144 16980 2148
rect 16996 2204 17060 2208
rect 16996 2148 17000 2204
rect 17000 2148 17056 2204
rect 17056 2148 17060 2204
rect 16996 2144 17060 2148
rect 17076 2204 17140 2208
rect 17076 2148 17080 2204
rect 17080 2148 17136 2204
rect 17136 2148 17140 2204
rect 17076 2144 17140 2148
rect 17156 2204 17220 2208
rect 17156 2148 17160 2204
rect 17160 2148 17216 2204
rect 17216 2148 17220 2204
rect 17156 2144 17220 2148
rect 17236 2204 17300 2208
rect 17236 2148 17240 2204
rect 17240 2148 17296 2204
rect 17296 2148 17300 2204
rect 17236 2144 17300 2148
rect 22916 2204 22980 2208
rect 22916 2148 22920 2204
rect 22920 2148 22976 2204
rect 22976 2148 22980 2204
rect 22916 2144 22980 2148
rect 22996 2204 23060 2208
rect 22996 2148 23000 2204
rect 23000 2148 23056 2204
rect 23056 2148 23060 2204
rect 22996 2144 23060 2148
rect 23076 2204 23140 2208
rect 23076 2148 23080 2204
rect 23080 2148 23136 2204
rect 23136 2148 23140 2204
rect 23076 2144 23140 2148
rect 23156 2204 23220 2208
rect 23156 2148 23160 2204
rect 23160 2148 23216 2204
rect 23216 2148 23220 2204
rect 23156 2144 23220 2148
rect 23236 2204 23300 2208
rect 23236 2148 23240 2204
rect 23240 2148 23296 2204
rect 23296 2148 23300 2204
rect 23236 2144 23300 2148
rect 28916 2204 28980 2208
rect 28916 2148 28920 2204
rect 28920 2148 28976 2204
rect 28976 2148 28980 2204
rect 28916 2144 28980 2148
rect 28996 2204 29060 2208
rect 28996 2148 29000 2204
rect 29000 2148 29056 2204
rect 29056 2148 29060 2204
rect 28996 2144 29060 2148
rect 29076 2204 29140 2208
rect 29076 2148 29080 2204
rect 29080 2148 29136 2204
rect 29136 2148 29140 2204
rect 29076 2144 29140 2148
rect 29156 2204 29220 2208
rect 29156 2148 29160 2204
rect 29160 2148 29216 2204
rect 29216 2148 29220 2204
rect 29156 2144 29220 2148
rect 29236 2204 29300 2208
rect 29236 2148 29240 2204
rect 29240 2148 29296 2204
rect 29296 2148 29300 2204
rect 29236 2144 29300 2148
<< metal4 >>
rect 4168 32128 4568 32144
rect 4168 32064 4176 32128
rect 4240 32064 4256 32128
rect 4320 32064 4336 32128
rect 4400 32064 4416 32128
rect 4480 32064 4496 32128
rect 4560 32064 4568 32128
rect 4168 31040 4568 32064
rect 4168 30976 4176 31040
rect 4240 30976 4256 31040
rect 4320 30976 4336 31040
rect 4400 30976 4416 31040
rect 4480 30976 4496 31040
rect 4560 30976 4568 31040
rect 4168 29952 4568 30976
rect 4168 29888 4176 29952
rect 4240 29888 4256 29952
rect 4320 29888 4336 29952
rect 4400 29888 4416 29952
rect 4480 29888 4496 29952
rect 4560 29888 4568 29952
rect 4168 29624 4568 29888
rect 4168 29388 4250 29624
rect 4486 29388 4568 29624
rect 4168 28864 4568 29388
rect 4168 28800 4176 28864
rect 4240 28800 4256 28864
rect 4320 28800 4336 28864
rect 4400 28800 4416 28864
rect 4480 28800 4496 28864
rect 4560 28800 4568 28864
rect 4168 27776 4568 28800
rect 4168 27712 4176 27776
rect 4240 27712 4256 27776
rect 4320 27712 4336 27776
rect 4400 27712 4416 27776
rect 4480 27712 4496 27776
rect 4560 27712 4568 27776
rect 4168 26688 4568 27712
rect 4168 26624 4176 26688
rect 4240 26624 4256 26688
rect 4320 26624 4336 26688
rect 4400 26624 4416 26688
rect 4480 26624 4496 26688
rect 4560 26624 4568 26688
rect 4168 25600 4568 26624
rect 4168 25536 4176 25600
rect 4240 25536 4256 25600
rect 4320 25536 4336 25600
rect 4400 25536 4416 25600
rect 4480 25536 4496 25600
rect 4560 25536 4568 25600
rect 4168 24512 4568 25536
rect 4168 24448 4176 24512
rect 4240 24448 4256 24512
rect 4320 24448 4336 24512
rect 4400 24448 4416 24512
rect 4480 24448 4496 24512
rect 4560 24448 4568 24512
rect 4168 23624 4568 24448
rect 4168 23424 4250 23624
rect 4486 23424 4568 23624
rect 4168 23360 4176 23424
rect 4240 23388 4250 23424
rect 4486 23388 4496 23424
rect 4240 23360 4256 23388
rect 4320 23360 4336 23388
rect 4400 23360 4416 23388
rect 4480 23360 4496 23388
rect 4560 23360 4568 23424
rect 4168 22336 4568 23360
rect 4168 22272 4176 22336
rect 4240 22272 4256 22336
rect 4320 22272 4336 22336
rect 4400 22272 4416 22336
rect 4480 22272 4496 22336
rect 4560 22272 4568 22336
rect 4168 21248 4568 22272
rect 4168 21184 4176 21248
rect 4240 21184 4256 21248
rect 4320 21184 4336 21248
rect 4400 21184 4416 21248
rect 4480 21184 4496 21248
rect 4560 21184 4568 21248
rect 4168 20160 4568 21184
rect 4168 20096 4176 20160
rect 4240 20096 4256 20160
rect 4320 20096 4336 20160
rect 4400 20096 4416 20160
rect 4480 20096 4496 20160
rect 4560 20096 4568 20160
rect 4168 19072 4568 20096
rect 4168 19008 4176 19072
rect 4240 19008 4256 19072
rect 4320 19008 4336 19072
rect 4400 19008 4416 19072
rect 4480 19008 4496 19072
rect 4560 19008 4568 19072
rect 4168 17984 4568 19008
rect 4168 17920 4176 17984
rect 4240 17920 4256 17984
rect 4320 17920 4336 17984
rect 4400 17920 4416 17984
rect 4480 17920 4496 17984
rect 4560 17920 4568 17984
rect 4168 17624 4568 17920
rect 4168 17388 4250 17624
rect 4486 17388 4568 17624
rect 4168 16896 4568 17388
rect 4168 16832 4176 16896
rect 4240 16832 4256 16896
rect 4320 16832 4336 16896
rect 4400 16832 4416 16896
rect 4480 16832 4496 16896
rect 4560 16832 4568 16896
rect 4168 15808 4568 16832
rect 4168 15744 4176 15808
rect 4240 15744 4256 15808
rect 4320 15744 4336 15808
rect 4400 15744 4416 15808
rect 4480 15744 4496 15808
rect 4560 15744 4568 15808
rect 4168 14720 4568 15744
rect 4168 14656 4176 14720
rect 4240 14656 4256 14720
rect 4320 14656 4336 14720
rect 4400 14656 4416 14720
rect 4480 14656 4496 14720
rect 4560 14656 4568 14720
rect 4168 13632 4568 14656
rect 4168 13568 4176 13632
rect 4240 13568 4256 13632
rect 4320 13568 4336 13632
rect 4400 13568 4416 13632
rect 4480 13568 4496 13632
rect 4560 13568 4568 13632
rect 4168 12544 4568 13568
rect 4168 12480 4176 12544
rect 4240 12480 4256 12544
rect 4320 12480 4336 12544
rect 4400 12480 4416 12544
rect 4480 12480 4496 12544
rect 4560 12480 4568 12544
rect 4168 11624 4568 12480
rect 4168 11456 4250 11624
rect 4486 11456 4568 11624
rect 4168 11392 4176 11456
rect 4240 11392 4250 11456
rect 4486 11392 4496 11456
rect 4560 11392 4568 11456
rect 4168 11388 4250 11392
rect 4486 11388 4568 11392
rect 4168 10368 4568 11388
rect 4168 10304 4176 10368
rect 4240 10304 4256 10368
rect 4320 10304 4336 10368
rect 4400 10304 4416 10368
rect 4480 10304 4496 10368
rect 4560 10304 4568 10368
rect 4168 9280 4568 10304
rect 4168 9216 4176 9280
rect 4240 9216 4256 9280
rect 4320 9216 4336 9280
rect 4400 9216 4416 9280
rect 4480 9216 4496 9280
rect 4560 9216 4568 9280
rect 4168 8192 4568 9216
rect 4168 8128 4176 8192
rect 4240 8128 4256 8192
rect 4320 8128 4336 8192
rect 4400 8128 4416 8192
rect 4480 8128 4496 8192
rect 4560 8128 4568 8192
rect 4168 7104 4568 8128
rect 4168 7040 4176 7104
rect 4240 7040 4256 7104
rect 4320 7040 4336 7104
rect 4400 7040 4416 7104
rect 4480 7040 4496 7104
rect 4560 7040 4568 7104
rect 4168 6016 4568 7040
rect 4168 5952 4176 6016
rect 4240 5952 4256 6016
rect 4320 5952 4336 6016
rect 4400 5952 4416 6016
rect 4480 5952 4496 6016
rect 4560 5952 4568 6016
rect 4168 5624 4568 5952
rect 4168 5388 4250 5624
rect 4486 5388 4568 5624
rect 4168 4928 4568 5388
rect 4168 4864 4176 4928
rect 4240 4864 4256 4928
rect 4320 4864 4336 4928
rect 4400 4864 4416 4928
rect 4480 4864 4496 4928
rect 4560 4864 4568 4928
rect 4168 3840 4568 4864
rect 4168 3776 4176 3840
rect 4240 3776 4256 3840
rect 4320 3776 4336 3840
rect 4400 3776 4416 3840
rect 4480 3776 4496 3840
rect 4560 3776 4568 3840
rect 4168 2752 4568 3776
rect 4168 2688 4176 2752
rect 4240 2688 4256 2752
rect 4320 2688 4336 2752
rect 4400 2688 4416 2752
rect 4480 2688 4496 2752
rect 4560 2688 4568 2752
rect 4168 2128 4568 2688
rect 4908 31584 5308 32144
rect 4908 31520 4916 31584
rect 4980 31520 4996 31584
rect 5060 31520 5076 31584
rect 5140 31520 5156 31584
rect 5220 31520 5236 31584
rect 5300 31520 5308 31584
rect 4908 30496 5308 31520
rect 4908 30432 4916 30496
rect 4980 30432 4996 30496
rect 5060 30432 5076 30496
rect 5140 30432 5156 30496
rect 5220 30432 5236 30496
rect 5300 30432 5308 30496
rect 4908 30364 5308 30432
rect 4908 30128 4990 30364
rect 5226 30128 5308 30364
rect 4908 29408 5308 30128
rect 4908 29344 4916 29408
rect 4980 29344 4996 29408
rect 5060 29344 5076 29408
rect 5140 29344 5156 29408
rect 5220 29344 5236 29408
rect 5300 29344 5308 29408
rect 4908 28320 5308 29344
rect 4908 28256 4916 28320
rect 4980 28256 4996 28320
rect 5060 28256 5076 28320
rect 5140 28256 5156 28320
rect 5220 28256 5236 28320
rect 5300 28256 5308 28320
rect 4908 27232 5308 28256
rect 4908 27168 4916 27232
rect 4980 27168 4996 27232
rect 5060 27168 5076 27232
rect 5140 27168 5156 27232
rect 5220 27168 5236 27232
rect 5300 27168 5308 27232
rect 4908 26144 5308 27168
rect 4908 26080 4916 26144
rect 4980 26080 4996 26144
rect 5060 26080 5076 26144
rect 5140 26080 5156 26144
rect 5220 26080 5236 26144
rect 5300 26080 5308 26144
rect 4908 25056 5308 26080
rect 4908 24992 4916 25056
rect 4980 24992 4996 25056
rect 5060 24992 5076 25056
rect 5140 24992 5156 25056
rect 5220 24992 5236 25056
rect 5300 24992 5308 25056
rect 4908 24364 5308 24992
rect 4908 24128 4990 24364
rect 5226 24128 5308 24364
rect 4908 23968 5308 24128
rect 4908 23904 4916 23968
rect 4980 23904 4996 23968
rect 5060 23904 5076 23968
rect 5140 23904 5156 23968
rect 5220 23904 5236 23968
rect 5300 23904 5308 23968
rect 4908 22880 5308 23904
rect 4908 22816 4916 22880
rect 4980 22816 4996 22880
rect 5060 22816 5076 22880
rect 5140 22816 5156 22880
rect 5220 22816 5236 22880
rect 5300 22816 5308 22880
rect 4908 21792 5308 22816
rect 4908 21728 4916 21792
rect 4980 21728 4996 21792
rect 5060 21728 5076 21792
rect 5140 21728 5156 21792
rect 5220 21728 5236 21792
rect 5300 21728 5308 21792
rect 4908 20704 5308 21728
rect 4908 20640 4916 20704
rect 4980 20640 4996 20704
rect 5060 20640 5076 20704
rect 5140 20640 5156 20704
rect 5220 20640 5236 20704
rect 5300 20640 5308 20704
rect 4908 19616 5308 20640
rect 4908 19552 4916 19616
rect 4980 19552 4996 19616
rect 5060 19552 5076 19616
rect 5140 19552 5156 19616
rect 5220 19552 5236 19616
rect 5300 19552 5308 19616
rect 4908 18528 5308 19552
rect 4908 18464 4916 18528
rect 4980 18464 4996 18528
rect 5060 18464 5076 18528
rect 5140 18464 5156 18528
rect 5220 18464 5236 18528
rect 5300 18464 5308 18528
rect 4908 18364 5308 18464
rect 4908 18128 4990 18364
rect 5226 18128 5308 18364
rect 4908 17440 5308 18128
rect 4908 17376 4916 17440
rect 4980 17376 4996 17440
rect 5060 17376 5076 17440
rect 5140 17376 5156 17440
rect 5220 17376 5236 17440
rect 5300 17376 5308 17440
rect 4908 16352 5308 17376
rect 4908 16288 4916 16352
rect 4980 16288 4996 16352
rect 5060 16288 5076 16352
rect 5140 16288 5156 16352
rect 5220 16288 5236 16352
rect 5300 16288 5308 16352
rect 4908 15264 5308 16288
rect 4908 15200 4916 15264
rect 4980 15200 4996 15264
rect 5060 15200 5076 15264
rect 5140 15200 5156 15264
rect 5220 15200 5236 15264
rect 5300 15200 5308 15264
rect 4908 14176 5308 15200
rect 4908 14112 4916 14176
rect 4980 14112 4996 14176
rect 5060 14112 5076 14176
rect 5140 14112 5156 14176
rect 5220 14112 5236 14176
rect 5300 14112 5308 14176
rect 4908 13088 5308 14112
rect 4908 13024 4916 13088
rect 4980 13024 4996 13088
rect 5060 13024 5076 13088
rect 5140 13024 5156 13088
rect 5220 13024 5236 13088
rect 5300 13024 5308 13088
rect 4908 12364 5308 13024
rect 4908 12128 4990 12364
rect 5226 12128 5308 12364
rect 4908 12000 5308 12128
rect 4908 11936 4916 12000
rect 4980 11936 4996 12000
rect 5060 11936 5076 12000
rect 5140 11936 5156 12000
rect 5220 11936 5236 12000
rect 5300 11936 5308 12000
rect 4908 10912 5308 11936
rect 4908 10848 4916 10912
rect 4980 10848 4996 10912
rect 5060 10848 5076 10912
rect 5140 10848 5156 10912
rect 5220 10848 5236 10912
rect 5300 10848 5308 10912
rect 4908 9824 5308 10848
rect 4908 9760 4916 9824
rect 4980 9760 4996 9824
rect 5060 9760 5076 9824
rect 5140 9760 5156 9824
rect 5220 9760 5236 9824
rect 5300 9760 5308 9824
rect 4908 8736 5308 9760
rect 4908 8672 4916 8736
rect 4980 8672 4996 8736
rect 5060 8672 5076 8736
rect 5140 8672 5156 8736
rect 5220 8672 5236 8736
rect 5300 8672 5308 8736
rect 4908 7648 5308 8672
rect 4908 7584 4916 7648
rect 4980 7584 4996 7648
rect 5060 7584 5076 7648
rect 5140 7584 5156 7648
rect 5220 7584 5236 7648
rect 5300 7584 5308 7648
rect 4908 6560 5308 7584
rect 4908 6496 4916 6560
rect 4980 6496 4996 6560
rect 5060 6496 5076 6560
rect 5140 6496 5156 6560
rect 5220 6496 5236 6560
rect 5300 6496 5308 6560
rect 4908 6364 5308 6496
rect 4908 6128 4990 6364
rect 5226 6128 5308 6364
rect 4908 5472 5308 6128
rect 4908 5408 4916 5472
rect 4980 5408 4996 5472
rect 5060 5408 5076 5472
rect 5140 5408 5156 5472
rect 5220 5408 5236 5472
rect 5300 5408 5308 5472
rect 4908 4384 5308 5408
rect 4908 4320 4916 4384
rect 4980 4320 4996 4384
rect 5060 4320 5076 4384
rect 5140 4320 5156 4384
rect 5220 4320 5236 4384
rect 5300 4320 5308 4384
rect 4908 3296 5308 4320
rect 4908 3232 4916 3296
rect 4980 3232 4996 3296
rect 5060 3232 5076 3296
rect 5140 3232 5156 3296
rect 5220 3232 5236 3296
rect 5300 3232 5308 3296
rect 4908 2208 5308 3232
rect 4908 2144 4916 2208
rect 4980 2144 4996 2208
rect 5060 2144 5076 2208
rect 5140 2144 5156 2208
rect 5220 2144 5236 2208
rect 5300 2144 5308 2208
rect 4908 2128 5308 2144
rect 10168 32128 10568 32144
rect 10168 32064 10176 32128
rect 10240 32064 10256 32128
rect 10320 32064 10336 32128
rect 10400 32064 10416 32128
rect 10480 32064 10496 32128
rect 10560 32064 10568 32128
rect 10168 31040 10568 32064
rect 10168 30976 10176 31040
rect 10240 30976 10256 31040
rect 10320 30976 10336 31040
rect 10400 30976 10416 31040
rect 10480 30976 10496 31040
rect 10560 30976 10568 31040
rect 10168 29952 10568 30976
rect 10168 29888 10176 29952
rect 10240 29888 10256 29952
rect 10320 29888 10336 29952
rect 10400 29888 10416 29952
rect 10480 29888 10496 29952
rect 10560 29888 10568 29952
rect 10168 29624 10568 29888
rect 10168 29388 10250 29624
rect 10486 29388 10568 29624
rect 10168 28864 10568 29388
rect 10168 28800 10176 28864
rect 10240 28800 10256 28864
rect 10320 28800 10336 28864
rect 10400 28800 10416 28864
rect 10480 28800 10496 28864
rect 10560 28800 10568 28864
rect 10168 27776 10568 28800
rect 10168 27712 10176 27776
rect 10240 27712 10256 27776
rect 10320 27712 10336 27776
rect 10400 27712 10416 27776
rect 10480 27712 10496 27776
rect 10560 27712 10568 27776
rect 10168 26688 10568 27712
rect 10168 26624 10176 26688
rect 10240 26624 10256 26688
rect 10320 26624 10336 26688
rect 10400 26624 10416 26688
rect 10480 26624 10496 26688
rect 10560 26624 10568 26688
rect 10168 25600 10568 26624
rect 10168 25536 10176 25600
rect 10240 25536 10256 25600
rect 10320 25536 10336 25600
rect 10400 25536 10416 25600
rect 10480 25536 10496 25600
rect 10560 25536 10568 25600
rect 10168 24512 10568 25536
rect 10168 24448 10176 24512
rect 10240 24448 10256 24512
rect 10320 24448 10336 24512
rect 10400 24448 10416 24512
rect 10480 24448 10496 24512
rect 10560 24448 10568 24512
rect 10168 23624 10568 24448
rect 10168 23424 10250 23624
rect 10486 23424 10568 23624
rect 10168 23360 10176 23424
rect 10240 23388 10250 23424
rect 10486 23388 10496 23424
rect 10240 23360 10256 23388
rect 10320 23360 10336 23388
rect 10400 23360 10416 23388
rect 10480 23360 10496 23388
rect 10560 23360 10568 23424
rect 10168 22336 10568 23360
rect 10168 22272 10176 22336
rect 10240 22272 10256 22336
rect 10320 22272 10336 22336
rect 10400 22272 10416 22336
rect 10480 22272 10496 22336
rect 10560 22272 10568 22336
rect 10168 21248 10568 22272
rect 10168 21184 10176 21248
rect 10240 21184 10256 21248
rect 10320 21184 10336 21248
rect 10400 21184 10416 21248
rect 10480 21184 10496 21248
rect 10560 21184 10568 21248
rect 10168 20160 10568 21184
rect 10168 20096 10176 20160
rect 10240 20096 10256 20160
rect 10320 20096 10336 20160
rect 10400 20096 10416 20160
rect 10480 20096 10496 20160
rect 10560 20096 10568 20160
rect 10168 19072 10568 20096
rect 10168 19008 10176 19072
rect 10240 19008 10256 19072
rect 10320 19008 10336 19072
rect 10400 19008 10416 19072
rect 10480 19008 10496 19072
rect 10560 19008 10568 19072
rect 10168 17984 10568 19008
rect 10168 17920 10176 17984
rect 10240 17920 10256 17984
rect 10320 17920 10336 17984
rect 10400 17920 10416 17984
rect 10480 17920 10496 17984
rect 10560 17920 10568 17984
rect 10168 17624 10568 17920
rect 10168 17388 10250 17624
rect 10486 17388 10568 17624
rect 10168 16896 10568 17388
rect 10168 16832 10176 16896
rect 10240 16832 10256 16896
rect 10320 16832 10336 16896
rect 10400 16832 10416 16896
rect 10480 16832 10496 16896
rect 10560 16832 10568 16896
rect 10168 15808 10568 16832
rect 10168 15744 10176 15808
rect 10240 15744 10256 15808
rect 10320 15744 10336 15808
rect 10400 15744 10416 15808
rect 10480 15744 10496 15808
rect 10560 15744 10568 15808
rect 10168 14720 10568 15744
rect 10168 14656 10176 14720
rect 10240 14656 10256 14720
rect 10320 14656 10336 14720
rect 10400 14656 10416 14720
rect 10480 14656 10496 14720
rect 10560 14656 10568 14720
rect 10168 13632 10568 14656
rect 10168 13568 10176 13632
rect 10240 13568 10256 13632
rect 10320 13568 10336 13632
rect 10400 13568 10416 13632
rect 10480 13568 10496 13632
rect 10560 13568 10568 13632
rect 10168 12544 10568 13568
rect 10168 12480 10176 12544
rect 10240 12480 10256 12544
rect 10320 12480 10336 12544
rect 10400 12480 10416 12544
rect 10480 12480 10496 12544
rect 10560 12480 10568 12544
rect 10168 11624 10568 12480
rect 10168 11456 10250 11624
rect 10486 11456 10568 11624
rect 10168 11392 10176 11456
rect 10240 11392 10250 11456
rect 10486 11392 10496 11456
rect 10560 11392 10568 11456
rect 10168 11388 10250 11392
rect 10486 11388 10568 11392
rect 10168 10368 10568 11388
rect 10168 10304 10176 10368
rect 10240 10304 10256 10368
rect 10320 10304 10336 10368
rect 10400 10304 10416 10368
rect 10480 10304 10496 10368
rect 10560 10304 10568 10368
rect 10168 9280 10568 10304
rect 10168 9216 10176 9280
rect 10240 9216 10256 9280
rect 10320 9216 10336 9280
rect 10400 9216 10416 9280
rect 10480 9216 10496 9280
rect 10560 9216 10568 9280
rect 10168 8192 10568 9216
rect 10168 8128 10176 8192
rect 10240 8128 10256 8192
rect 10320 8128 10336 8192
rect 10400 8128 10416 8192
rect 10480 8128 10496 8192
rect 10560 8128 10568 8192
rect 10168 7104 10568 8128
rect 10168 7040 10176 7104
rect 10240 7040 10256 7104
rect 10320 7040 10336 7104
rect 10400 7040 10416 7104
rect 10480 7040 10496 7104
rect 10560 7040 10568 7104
rect 10168 6016 10568 7040
rect 10168 5952 10176 6016
rect 10240 5952 10256 6016
rect 10320 5952 10336 6016
rect 10400 5952 10416 6016
rect 10480 5952 10496 6016
rect 10560 5952 10568 6016
rect 10168 5624 10568 5952
rect 10168 5388 10250 5624
rect 10486 5388 10568 5624
rect 10168 4928 10568 5388
rect 10168 4864 10176 4928
rect 10240 4864 10256 4928
rect 10320 4864 10336 4928
rect 10400 4864 10416 4928
rect 10480 4864 10496 4928
rect 10560 4864 10568 4928
rect 10168 3840 10568 4864
rect 10168 3776 10176 3840
rect 10240 3776 10256 3840
rect 10320 3776 10336 3840
rect 10400 3776 10416 3840
rect 10480 3776 10496 3840
rect 10560 3776 10568 3840
rect 10168 2752 10568 3776
rect 10168 2688 10176 2752
rect 10240 2688 10256 2752
rect 10320 2688 10336 2752
rect 10400 2688 10416 2752
rect 10480 2688 10496 2752
rect 10560 2688 10568 2752
rect 10168 2128 10568 2688
rect 10908 31584 11308 32144
rect 10908 31520 10916 31584
rect 10980 31520 10996 31584
rect 11060 31520 11076 31584
rect 11140 31520 11156 31584
rect 11220 31520 11236 31584
rect 11300 31520 11308 31584
rect 10908 30496 11308 31520
rect 10908 30432 10916 30496
rect 10980 30432 10996 30496
rect 11060 30432 11076 30496
rect 11140 30432 11156 30496
rect 11220 30432 11236 30496
rect 11300 30432 11308 30496
rect 10908 30364 11308 30432
rect 10908 30128 10990 30364
rect 11226 30128 11308 30364
rect 10908 29408 11308 30128
rect 10908 29344 10916 29408
rect 10980 29344 10996 29408
rect 11060 29344 11076 29408
rect 11140 29344 11156 29408
rect 11220 29344 11236 29408
rect 11300 29344 11308 29408
rect 10908 28320 11308 29344
rect 10908 28256 10916 28320
rect 10980 28256 10996 28320
rect 11060 28256 11076 28320
rect 11140 28256 11156 28320
rect 11220 28256 11236 28320
rect 11300 28256 11308 28320
rect 10908 27232 11308 28256
rect 10908 27168 10916 27232
rect 10980 27168 10996 27232
rect 11060 27168 11076 27232
rect 11140 27168 11156 27232
rect 11220 27168 11236 27232
rect 11300 27168 11308 27232
rect 10908 26144 11308 27168
rect 10908 26080 10916 26144
rect 10980 26080 10996 26144
rect 11060 26080 11076 26144
rect 11140 26080 11156 26144
rect 11220 26080 11236 26144
rect 11300 26080 11308 26144
rect 10908 25056 11308 26080
rect 10908 24992 10916 25056
rect 10980 24992 10996 25056
rect 11060 24992 11076 25056
rect 11140 24992 11156 25056
rect 11220 24992 11236 25056
rect 11300 24992 11308 25056
rect 10908 24364 11308 24992
rect 10908 24128 10990 24364
rect 11226 24128 11308 24364
rect 10908 23968 11308 24128
rect 10908 23904 10916 23968
rect 10980 23904 10996 23968
rect 11060 23904 11076 23968
rect 11140 23904 11156 23968
rect 11220 23904 11236 23968
rect 11300 23904 11308 23968
rect 10908 22880 11308 23904
rect 16168 32128 16568 32144
rect 16168 32064 16176 32128
rect 16240 32064 16256 32128
rect 16320 32064 16336 32128
rect 16400 32064 16416 32128
rect 16480 32064 16496 32128
rect 16560 32064 16568 32128
rect 16168 31040 16568 32064
rect 16168 30976 16176 31040
rect 16240 30976 16256 31040
rect 16320 30976 16336 31040
rect 16400 30976 16416 31040
rect 16480 30976 16496 31040
rect 16560 30976 16568 31040
rect 16168 29952 16568 30976
rect 16168 29888 16176 29952
rect 16240 29888 16256 29952
rect 16320 29888 16336 29952
rect 16400 29888 16416 29952
rect 16480 29888 16496 29952
rect 16560 29888 16568 29952
rect 16168 29624 16568 29888
rect 16168 29388 16250 29624
rect 16486 29388 16568 29624
rect 16168 28864 16568 29388
rect 16168 28800 16176 28864
rect 16240 28800 16256 28864
rect 16320 28800 16336 28864
rect 16400 28800 16416 28864
rect 16480 28800 16496 28864
rect 16560 28800 16568 28864
rect 16168 27776 16568 28800
rect 16168 27712 16176 27776
rect 16240 27712 16256 27776
rect 16320 27712 16336 27776
rect 16400 27712 16416 27776
rect 16480 27712 16496 27776
rect 16560 27712 16568 27776
rect 16168 26688 16568 27712
rect 16168 26624 16176 26688
rect 16240 26624 16256 26688
rect 16320 26624 16336 26688
rect 16400 26624 16416 26688
rect 16480 26624 16496 26688
rect 16560 26624 16568 26688
rect 16168 25600 16568 26624
rect 16168 25536 16176 25600
rect 16240 25536 16256 25600
rect 16320 25536 16336 25600
rect 16400 25536 16416 25600
rect 16480 25536 16496 25600
rect 16560 25536 16568 25600
rect 16168 24512 16568 25536
rect 16168 24448 16176 24512
rect 16240 24448 16256 24512
rect 16320 24448 16336 24512
rect 16400 24448 16416 24512
rect 16480 24448 16496 24512
rect 16560 24448 16568 24512
rect 15331 23628 15397 23629
rect 15331 23564 15332 23628
rect 15396 23564 15397 23628
rect 15331 23563 15397 23564
rect 16168 23624 16568 24448
rect 10908 22816 10916 22880
rect 10980 22816 10996 22880
rect 11060 22816 11076 22880
rect 11140 22816 11156 22880
rect 11220 22816 11236 22880
rect 11300 22816 11308 22880
rect 10908 21792 11308 22816
rect 10908 21728 10916 21792
rect 10980 21728 10996 21792
rect 11060 21728 11076 21792
rect 11140 21728 11156 21792
rect 11220 21728 11236 21792
rect 11300 21728 11308 21792
rect 10908 20704 11308 21728
rect 10908 20640 10916 20704
rect 10980 20640 10996 20704
rect 11060 20640 11076 20704
rect 11140 20640 11156 20704
rect 11220 20640 11236 20704
rect 11300 20640 11308 20704
rect 10908 19616 11308 20640
rect 10908 19552 10916 19616
rect 10980 19552 10996 19616
rect 11060 19552 11076 19616
rect 11140 19552 11156 19616
rect 11220 19552 11236 19616
rect 11300 19552 11308 19616
rect 10908 18528 11308 19552
rect 10908 18464 10916 18528
rect 10980 18464 10996 18528
rect 11060 18464 11076 18528
rect 11140 18464 11156 18528
rect 11220 18464 11236 18528
rect 11300 18464 11308 18528
rect 10908 18364 11308 18464
rect 10908 18128 10990 18364
rect 11226 18128 11308 18364
rect 10908 17440 11308 18128
rect 10908 17376 10916 17440
rect 10980 17376 10996 17440
rect 11060 17376 11076 17440
rect 11140 17376 11156 17440
rect 11220 17376 11236 17440
rect 11300 17376 11308 17440
rect 10908 16352 11308 17376
rect 15334 17373 15394 23563
rect 16168 23424 16250 23624
rect 16486 23424 16568 23624
rect 16168 23360 16176 23424
rect 16240 23388 16250 23424
rect 16486 23388 16496 23424
rect 16240 23360 16256 23388
rect 16320 23360 16336 23388
rect 16400 23360 16416 23388
rect 16480 23360 16496 23388
rect 16560 23360 16568 23424
rect 16168 22336 16568 23360
rect 16168 22272 16176 22336
rect 16240 22272 16256 22336
rect 16320 22272 16336 22336
rect 16400 22272 16416 22336
rect 16480 22272 16496 22336
rect 16560 22272 16568 22336
rect 16168 21248 16568 22272
rect 16168 21184 16176 21248
rect 16240 21184 16256 21248
rect 16320 21184 16336 21248
rect 16400 21184 16416 21248
rect 16480 21184 16496 21248
rect 16560 21184 16568 21248
rect 16168 20160 16568 21184
rect 16168 20096 16176 20160
rect 16240 20096 16256 20160
rect 16320 20096 16336 20160
rect 16400 20096 16416 20160
rect 16480 20096 16496 20160
rect 16560 20096 16568 20160
rect 16168 19072 16568 20096
rect 16168 19008 16176 19072
rect 16240 19008 16256 19072
rect 16320 19008 16336 19072
rect 16400 19008 16416 19072
rect 16480 19008 16496 19072
rect 16560 19008 16568 19072
rect 16168 17984 16568 19008
rect 16168 17920 16176 17984
rect 16240 17920 16256 17984
rect 16320 17920 16336 17984
rect 16400 17920 16416 17984
rect 16480 17920 16496 17984
rect 16560 17920 16568 17984
rect 16168 17624 16568 17920
rect 16168 17388 16250 17624
rect 16486 17388 16568 17624
rect 15331 17372 15397 17373
rect 15331 17308 15332 17372
rect 15396 17308 15397 17372
rect 15331 17307 15397 17308
rect 10908 16288 10916 16352
rect 10980 16288 10996 16352
rect 11060 16288 11076 16352
rect 11140 16288 11156 16352
rect 11220 16288 11236 16352
rect 11300 16288 11308 16352
rect 10908 15264 11308 16288
rect 10908 15200 10916 15264
rect 10980 15200 10996 15264
rect 11060 15200 11076 15264
rect 11140 15200 11156 15264
rect 11220 15200 11236 15264
rect 11300 15200 11308 15264
rect 10908 14176 11308 15200
rect 10908 14112 10916 14176
rect 10980 14112 10996 14176
rect 11060 14112 11076 14176
rect 11140 14112 11156 14176
rect 11220 14112 11236 14176
rect 11300 14112 11308 14176
rect 10908 13088 11308 14112
rect 10908 13024 10916 13088
rect 10980 13024 10996 13088
rect 11060 13024 11076 13088
rect 11140 13024 11156 13088
rect 11220 13024 11236 13088
rect 11300 13024 11308 13088
rect 10908 12364 11308 13024
rect 15334 12885 15394 17307
rect 16168 16896 16568 17388
rect 16168 16832 16176 16896
rect 16240 16832 16256 16896
rect 16320 16832 16336 16896
rect 16400 16832 16416 16896
rect 16480 16832 16496 16896
rect 16560 16832 16568 16896
rect 16168 15808 16568 16832
rect 16168 15744 16176 15808
rect 16240 15744 16256 15808
rect 16320 15744 16336 15808
rect 16400 15744 16416 15808
rect 16480 15744 16496 15808
rect 16560 15744 16568 15808
rect 16168 14720 16568 15744
rect 16168 14656 16176 14720
rect 16240 14656 16256 14720
rect 16320 14656 16336 14720
rect 16400 14656 16416 14720
rect 16480 14656 16496 14720
rect 16560 14656 16568 14720
rect 16168 13632 16568 14656
rect 16168 13568 16176 13632
rect 16240 13568 16256 13632
rect 16320 13568 16336 13632
rect 16400 13568 16416 13632
rect 16480 13568 16496 13632
rect 16560 13568 16568 13632
rect 15331 12884 15397 12885
rect 15331 12820 15332 12884
rect 15396 12820 15397 12884
rect 15331 12819 15397 12820
rect 10908 12128 10990 12364
rect 11226 12128 11308 12364
rect 10908 12000 11308 12128
rect 10908 11936 10916 12000
rect 10980 11936 10996 12000
rect 11060 11936 11076 12000
rect 11140 11936 11156 12000
rect 11220 11936 11236 12000
rect 11300 11936 11308 12000
rect 10908 10912 11308 11936
rect 15334 11117 15394 12819
rect 16168 12544 16568 13568
rect 16168 12480 16176 12544
rect 16240 12480 16256 12544
rect 16320 12480 16336 12544
rect 16400 12480 16416 12544
rect 16480 12480 16496 12544
rect 16560 12480 16568 12544
rect 16168 11624 16568 12480
rect 16168 11456 16250 11624
rect 16486 11456 16568 11624
rect 16168 11392 16176 11456
rect 16240 11392 16250 11456
rect 16486 11392 16496 11456
rect 16560 11392 16568 11456
rect 16168 11388 16250 11392
rect 16486 11388 16568 11392
rect 15331 11116 15397 11117
rect 15331 11052 15332 11116
rect 15396 11052 15397 11116
rect 15331 11051 15397 11052
rect 10908 10848 10916 10912
rect 10980 10848 10996 10912
rect 11060 10848 11076 10912
rect 11140 10848 11156 10912
rect 11220 10848 11236 10912
rect 11300 10848 11308 10912
rect 10908 9824 11308 10848
rect 10908 9760 10916 9824
rect 10980 9760 10996 9824
rect 11060 9760 11076 9824
rect 11140 9760 11156 9824
rect 11220 9760 11236 9824
rect 11300 9760 11308 9824
rect 10908 8736 11308 9760
rect 10908 8672 10916 8736
rect 10980 8672 10996 8736
rect 11060 8672 11076 8736
rect 11140 8672 11156 8736
rect 11220 8672 11236 8736
rect 11300 8672 11308 8736
rect 10908 7648 11308 8672
rect 10908 7584 10916 7648
rect 10980 7584 10996 7648
rect 11060 7584 11076 7648
rect 11140 7584 11156 7648
rect 11220 7584 11236 7648
rect 11300 7584 11308 7648
rect 10908 6560 11308 7584
rect 10908 6496 10916 6560
rect 10980 6496 10996 6560
rect 11060 6496 11076 6560
rect 11140 6496 11156 6560
rect 11220 6496 11236 6560
rect 11300 6496 11308 6560
rect 10908 6364 11308 6496
rect 10908 6128 10990 6364
rect 11226 6128 11308 6364
rect 10908 5472 11308 6128
rect 10908 5408 10916 5472
rect 10980 5408 10996 5472
rect 11060 5408 11076 5472
rect 11140 5408 11156 5472
rect 11220 5408 11236 5472
rect 11300 5408 11308 5472
rect 10908 4384 11308 5408
rect 10908 4320 10916 4384
rect 10980 4320 10996 4384
rect 11060 4320 11076 4384
rect 11140 4320 11156 4384
rect 11220 4320 11236 4384
rect 11300 4320 11308 4384
rect 10908 3296 11308 4320
rect 10908 3232 10916 3296
rect 10980 3232 10996 3296
rect 11060 3232 11076 3296
rect 11140 3232 11156 3296
rect 11220 3232 11236 3296
rect 11300 3232 11308 3296
rect 10908 2208 11308 3232
rect 10908 2144 10916 2208
rect 10980 2144 10996 2208
rect 11060 2144 11076 2208
rect 11140 2144 11156 2208
rect 11220 2144 11236 2208
rect 11300 2144 11308 2208
rect 10908 2128 11308 2144
rect 16168 10368 16568 11388
rect 16168 10304 16176 10368
rect 16240 10304 16256 10368
rect 16320 10304 16336 10368
rect 16400 10304 16416 10368
rect 16480 10304 16496 10368
rect 16560 10304 16568 10368
rect 16168 9280 16568 10304
rect 16168 9216 16176 9280
rect 16240 9216 16256 9280
rect 16320 9216 16336 9280
rect 16400 9216 16416 9280
rect 16480 9216 16496 9280
rect 16560 9216 16568 9280
rect 16168 8192 16568 9216
rect 16168 8128 16176 8192
rect 16240 8128 16256 8192
rect 16320 8128 16336 8192
rect 16400 8128 16416 8192
rect 16480 8128 16496 8192
rect 16560 8128 16568 8192
rect 16168 7104 16568 8128
rect 16168 7040 16176 7104
rect 16240 7040 16256 7104
rect 16320 7040 16336 7104
rect 16400 7040 16416 7104
rect 16480 7040 16496 7104
rect 16560 7040 16568 7104
rect 16168 6016 16568 7040
rect 16168 5952 16176 6016
rect 16240 5952 16256 6016
rect 16320 5952 16336 6016
rect 16400 5952 16416 6016
rect 16480 5952 16496 6016
rect 16560 5952 16568 6016
rect 16168 5624 16568 5952
rect 16168 5388 16250 5624
rect 16486 5388 16568 5624
rect 16168 4928 16568 5388
rect 16168 4864 16176 4928
rect 16240 4864 16256 4928
rect 16320 4864 16336 4928
rect 16400 4864 16416 4928
rect 16480 4864 16496 4928
rect 16560 4864 16568 4928
rect 16168 3840 16568 4864
rect 16168 3776 16176 3840
rect 16240 3776 16256 3840
rect 16320 3776 16336 3840
rect 16400 3776 16416 3840
rect 16480 3776 16496 3840
rect 16560 3776 16568 3840
rect 16168 2752 16568 3776
rect 16168 2688 16176 2752
rect 16240 2688 16256 2752
rect 16320 2688 16336 2752
rect 16400 2688 16416 2752
rect 16480 2688 16496 2752
rect 16560 2688 16568 2752
rect 16168 2128 16568 2688
rect 16908 31584 17308 32144
rect 16908 31520 16916 31584
rect 16980 31520 16996 31584
rect 17060 31520 17076 31584
rect 17140 31520 17156 31584
rect 17220 31520 17236 31584
rect 17300 31520 17308 31584
rect 16908 30496 17308 31520
rect 16908 30432 16916 30496
rect 16980 30432 16996 30496
rect 17060 30432 17076 30496
rect 17140 30432 17156 30496
rect 17220 30432 17236 30496
rect 17300 30432 17308 30496
rect 16908 30364 17308 30432
rect 16908 30128 16990 30364
rect 17226 30128 17308 30364
rect 16908 29408 17308 30128
rect 16908 29344 16916 29408
rect 16980 29344 16996 29408
rect 17060 29344 17076 29408
rect 17140 29344 17156 29408
rect 17220 29344 17236 29408
rect 17300 29344 17308 29408
rect 16908 28320 17308 29344
rect 16908 28256 16916 28320
rect 16980 28256 16996 28320
rect 17060 28256 17076 28320
rect 17140 28256 17156 28320
rect 17220 28256 17236 28320
rect 17300 28256 17308 28320
rect 16908 27232 17308 28256
rect 16908 27168 16916 27232
rect 16980 27168 16996 27232
rect 17060 27168 17076 27232
rect 17140 27168 17156 27232
rect 17220 27168 17236 27232
rect 17300 27168 17308 27232
rect 16908 26144 17308 27168
rect 22168 32128 22568 32144
rect 22168 32064 22176 32128
rect 22240 32064 22256 32128
rect 22320 32064 22336 32128
rect 22400 32064 22416 32128
rect 22480 32064 22496 32128
rect 22560 32064 22568 32128
rect 22168 31040 22568 32064
rect 22168 30976 22176 31040
rect 22240 30976 22256 31040
rect 22320 30976 22336 31040
rect 22400 30976 22416 31040
rect 22480 30976 22496 31040
rect 22560 30976 22568 31040
rect 22168 29952 22568 30976
rect 22168 29888 22176 29952
rect 22240 29888 22256 29952
rect 22320 29888 22336 29952
rect 22400 29888 22416 29952
rect 22480 29888 22496 29952
rect 22560 29888 22568 29952
rect 22168 29624 22568 29888
rect 22168 29388 22250 29624
rect 22486 29388 22568 29624
rect 22168 28864 22568 29388
rect 22168 28800 22176 28864
rect 22240 28800 22256 28864
rect 22320 28800 22336 28864
rect 22400 28800 22416 28864
rect 22480 28800 22496 28864
rect 22560 28800 22568 28864
rect 22168 27776 22568 28800
rect 22168 27712 22176 27776
rect 22240 27712 22256 27776
rect 22320 27712 22336 27776
rect 22400 27712 22416 27776
rect 22480 27712 22496 27776
rect 22560 27712 22568 27776
rect 22168 26688 22568 27712
rect 22168 26624 22176 26688
rect 22240 26624 22256 26688
rect 22320 26624 22336 26688
rect 22400 26624 22416 26688
rect 22480 26624 22496 26688
rect 22560 26624 22568 26688
rect 18643 26348 18709 26349
rect 18643 26284 18644 26348
rect 18708 26284 18709 26348
rect 18643 26283 18709 26284
rect 16908 26080 16916 26144
rect 16980 26080 16996 26144
rect 17060 26080 17076 26144
rect 17140 26080 17156 26144
rect 17220 26080 17236 26144
rect 17300 26080 17308 26144
rect 16908 25056 17308 26080
rect 16908 24992 16916 25056
rect 16980 24992 16996 25056
rect 17060 24992 17076 25056
rect 17140 24992 17156 25056
rect 17220 24992 17236 25056
rect 17300 24992 17308 25056
rect 16908 24364 17308 24992
rect 16908 24128 16990 24364
rect 17226 24128 17308 24364
rect 16908 23968 17308 24128
rect 16908 23904 16916 23968
rect 16980 23904 16996 23968
rect 17060 23904 17076 23968
rect 17140 23904 17156 23968
rect 17220 23904 17236 23968
rect 17300 23904 17308 23968
rect 16908 22880 17308 23904
rect 16908 22816 16916 22880
rect 16980 22816 16996 22880
rect 17060 22816 17076 22880
rect 17140 22816 17156 22880
rect 17220 22816 17236 22880
rect 17300 22816 17308 22880
rect 16908 21792 17308 22816
rect 16908 21728 16916 21792
rect 16980 21728 16996 21792
rect 17060 21728 17076 21792
rect 17140 21728 17156 21792
rect 17220 21728 17236 21792
rect 17300 21728 17308 21792
rect 16908 20704 17308 21728
rect 16908 20640 16916 20704
rect 16980 20640 16996 20704
rect 17060 20640 17076 20704
rect 17140 20640 17156 20704
rect 17220 20640 17236 20704
rect 17300 20640 17308 20704
rect 16908 19616 17308 20640
rect 16908 19552 16916 19616
rect 16980 19552 16996 19616
rect 17060 19552 17076 19616
rect 17140 19552 17156 19616
rect 17220 19552 17236 19616
rect 17300 19552 17308 19616
rect 16908 18528 17308 19552
rect 16908 18464 16916 18528
rect 16980 18464 16996 18528
rect 17060 18464 17076 18528
rect 17140 18464 17156 18528
rect 17220 18464 17236 18528
rect 17300 18464 17308 18528
rect 16908 18364 17308 18464
rect 16908 18128 16990 18364
rect 17226 18128 17308 18364
rect 16908 17440 17308 18128
rect 16908 17376 16916 17440
rect 16980 17376 16996 17440
rect 17060 17376 17076 17440
rect 17140 17376 17156 17440
rect 17220 17376 17236 17440
rect 17300 17376 17308 17440
rect 16908 16352 17308 17376
rect 16908 16288 16916 16352
rect 16980 16288 16996 16352
rect 17060 16288 17076 16352
rect 17140 16288 17156 16352
rect 17220 16288 17236 16352
rect 17300 16288 17308 16352
rect 16908 15264 17308 16288
rect 16908 15200 16916 15264
rect 16980 15200 16996 15264
rect 17060 15200 17076 15264
rect 17140 15200 17156 15264
rect 17220 15200 17236 15264
rect 17300 15200 17308 15264
rect 16908 14176 17308 15200
rect 16908 14112 16916 14176
rect 16980 14112 16996 14176
rect 17060 14112 17076 14176
rect 17140 14112 17156 14176
rect 17220 14112 17236 14176
rect 17300 14112 17308 14176
rect 16908 13088 17308 14112
rect 16908 13024 16916 13088
rect 16980 13024 16996 13088
rect 17060 13024 17076 13088
rect 17140 13024 17156 13088
rect 17220 13024 17236 13088
rect 17300 13024 17308 13088
rect 16908 12364 17308 13024
rect 16908 12128 16990 12364
rect 17226 12128 17308 12364
rect 16908 12000 17308 12128
rect 16908 11936 16916 12000
rect 16980 11936 16996 12000
rect 17060 11936 17076 12000
rect 17140 11936 17156 12000
rect 17220 11936 17236 12000
rect 17300 11936 17308 12000
rect 16908 10912 17308 11936
rect 16908 10848 16916 10912
rect 16980 10848 16996 10912
rect 17060 10848 17076 10912
rect 17140 10848 17156 10912
rect 17220 10848 17236 10912
rect 17300 10848 17308 10912
rect 16908 9824 17308 10848
rect 16908 9760 16916 9824
rect 16980 9760 16996 9824
rect 17060 9760 17076 9824
rect 17140 9760 17156 9824
rect 17220 9760 17236 9824
rect 17300 9760 17308 9824
rect 16908 8736 17308 9760
rect 18646 8805 18706 26283
rect 22168 25600 22568 26624
rect 22168 25536 22176 25600
rect 22240 25536 22256 25600
rect 22320 25536 22336 25600
rect 22400 25536 22416 25600
rect 22480 25536 22496 25600
rect 22560 25536 22568 25600
rect 22168 24512 22568 25536
rect 22168 24448 22176 24512
rect 22240 24448 22256 24512
rect 22320 24448 22336 24512
rect 22400 24448 22416 24512
rect 22480 24448 22496 24512
rect 22560 24448 22568 24512
rect 22168 23624 22568 24448
rect 22168 23424 22250 23624
rect 22486 23424 22568 23624
rect 22168 23360 22176 23424
rect 22240 23388 22250 23424
rect 22486 23388 22496 23424
rect 22240 23360 22256 23388
rect 22320 23360 22336 23388
rect 22400 23360 22416 23388
rect 22480 23360 22496 23388
rect 22560 23360 22568 23424
rect 22168 22336 22568 23360
rect 22168 22272 22176 22336
rect 22240 22272 22256 22336
rect 22320 22272 22336 22336
rect 22400 22272 22416 22336
rect 22480 22272 22496 22336
rect 22560 22272 22568 22336
rect 22168 21248 22568 22272
rect 22168 21184 22176 21248
rect 22240 21184 22256 21248
rect 22320 21184 22336 21248
rect 22400 21184 22416 21248
rect 22480 21184 22496 21248
rect 22560 21184 22568 21248
rect 22168 20160 22568 21184
rect 22168 20096 22176 20160
rect 22240 20096 22256 20160
rect 22320 20096 22336 20160
rect 22400 20096 22416 20160
rect 22480 20096 22496 20160
rect 22560 20096 22568 20160
rect 22168 19072 22568 20096
rect 22168 19008 22176 19072
rect 22240 19008 22256 19072
rect 22320 19008 22336 19072
rect 22400 19008 22416 19072
rect 22480 19008 22496 19072
rect 22560 19008 22568 19072
rect 22168 17984 22568 19008
rect 22168 17920 22176 17984
rect 22240 17920 22256 17984
rect 22320 17920 22336 17984
rect 22400 17920 22416 17984
rect 22480 17920 22496 17984
rect 22560 17920 22568 17984
rect 22168 17624 22568 17920
rect 22168 17388 22250 17624
rect 22486 17388 22568 17624
rect 22168 16896 22568 17388
rect 22168 16832 22176 16896
rect 22240 16832 22256 16896
rect 22320 16832 22336 16896
rect 22400 16832 22416 16896
rect 22480 16832 22496 16896
rect 22560 16832 22568 16896
rect 22168 15808 22568 16832
rect 22168 15744 22176 15808
rect 22240 15744 22256 15808
rect 22320 15744 22336 15808
rect 22400 15744 22416 15808
rect 22480 15744 22496 15808
rect 22560 15744 22568 15808
rect 22168 14720 22568 15744
rect 22168 14656 22176 14720
rect 22240 14656 22256 14720
rect 22320 14656 22336 14720
rect 22400 14656 22416 14720
rect 22480 14656 22496 14720
rect 22560 14656 22568 14720
rect 22168 13632 22568 14656
rect 22168 13568 22176 13632
rect 22240 13568 22256 13632
rect 22320 13568 22336 13632
rect 22400 13568 22416 13632
rect 22480 13568 22496 13632
rect 22560 13568 22568 13632
rect 22168 12544 22568 13568
rect 22168 12480 22176 12544
rect 22240 12480 22256 12544
rect 22320 12480 22336 12544
rect 22400 12480 22416 12544
rect 22480 12480 22496 12544
rect 22560 12480 22568 12544
rect 22168 11624 22568 12480
rect 22168 11456 22250 11624
rect 22486 11456 22568 11624
rect 22168 11392 22176 11456
rect 22240 11392 22250 11456
rect 22486 11392 22496 11456
rect 22560 11392 22568 11456
rect 22168 11388 22250 11392
rect 22486 11388 22568 11392
rect 22168 10368 22568 11388
rect 22168 10304 22176 10368
rect 22240 10304 22256 10368
rect 22320 10304 22336 10368
rect 22400 10304 22416 10368
rect 22480 10304 22496 10368
rect 22560 10304 22568 10368
rect 22168 9280 22568 10304
rect 22168 9216 22176 9280
rect 22240 9216 22256 9280
rect 22320 9216 22336 9280
rect 22400 9216 22416 9280
rect 22480 9216 22496 9280
rect 22560 9216 22568 9280
rect 18643 8804 18709 8805
rect 18643 8740 18644 8804
rect 18708 8740 18709 8804
rect 18643 8739 18709 8740
rect 16908 8672 16916 8736
rect 16980 8672 16996 8736
rect 17060 8672 17076 8736
rect 17140 8672 17156 8736
rect 17220 8672 17236 8736
rect 17300 8672 17308 8736
rect 16908 7648 17308 8672
rect 16908 7584 16916 7648
rect 16980 7584 16996 7648
rect 17060 7584 17076 7648
rect 17140 7584 17156 7648
rect 17220 7584 17236 7648
rect 17300 7584 17308 7648
rect 16908 6560 17308 7584
rect 16908 6496 16916 6560
rect 16980 6496 16996 6560
rect 17060 6496 17076 6560
rect 17140 6496 17156 6560
rect 17220 6496 17236 6560
rect 17300 6496 17308 6560
rect 16908 6364 17308 6496
rect 16908 6128 16990 6364
rect 17226 6128 17308 6364
rect 16908 5472 17308 6128
rect 16908 5408 16916 5472
rect 16980 5408 16996 5472
rect 17060 5408 17076 5472
rect 17140 5408 17156 5472
rect 17220 5408 17236 5472
rect 17300 5408 17308 5472
rect 16908 4384 17308 5408
rect 16908 4320 16916 4384
rect 16980 4320 16996 4384
rect 17060 4320 17076 4384
rect 17140 4320 17156 4384
rect 17220 4320 17236 4384
rect 17300 4320 17308 4384
rect 16908 3296 17308 4320
rect 16908 3232 16916 3296
rect 16980 3232 16996 3296
rect 17060 3232 17076 3296
rect 17140 3232 17156 3296
rect 17220 3232 17236 3296
rect 17300 3232 17308 3296
rect 16908 2208 17308 3232
rect 16908 2144 16916 2208
rect 16980 2144 16996 2208
rect 17060 2144 17076 2208
rect 17140 2144 17156 2208
rect 17220 2144 17236 2208
rect 17300 2144 17308 2208
rect 16908 2128 17308 2144
rect 22168 8192 22568 9216
rect 22168 8128 22176 8192
rect 22240 8128 22256 8192
rect 22320 8128 22336 8192
rect 22400 8128 22416 8192
rect 22480 8128 22496 8192
rect 22560 8128 22568 8192
rect 22168 7104 22568 8128
rect 22168 7040 22176 7104
rect 22240 7040 22256 7104
rect 22320 7040 22336 7104
rect 22400 7040 22416 7104
rect 22480 7040 22496 7104
rect 22560 7040 22568 7104
rect 22168 6016 22568 7040
rect 22168 5952 22176 6016
rect 22240 5952 22256 6016
rect 22320 5952 22336 6016
rect 22400 5952 22416 6016
rect 22480 5952 22496 6016
rect 22560 5952 22568 6016
rect 22168 5624 22568 5952
rect 22168 5388 22250 5624
rect 22486 5388 22568 5624
rect 22168 4928 22568 5388
rect 22168 4864 22176 4928
rect 22240 4864 22256 4928
rect 22320 4864 22336 4928
rect 22400 4864 22416 4928
rect 22480 4864 22496 4928
rect 22560 4864 22568 4928
rect 22168 3840 22568 4864
rect 22168 3776 22176 3840
rect 22240 3776 22256 3840
rect 22320 3776 22336 3840
rect 22400 3776 22416 3840
rect 22480 3776 22496 3840
rect 22560 3776 22568 3840
rect 22168 2752 22568 3776
rect 22168 2688 22176 2752
rect 22240 2688 22256 2752
rect 22320 2688 22336 2752
rect 22400 2688 22416 2752
rect 22480 2688 22496 2752
rect 22560 2688 22568 2752
rect 22168 2128 22568 2688
rect 22908 31584 23308 32144
rect 28168 32128 28568 32144
rect 28168 32064 28176 32128
rect 28240 32064 28256 32128
rect 28320 32064 28336 32128
rect 28400 32064 28416 32128
rect 28480 32064 28496 32128
rect 28560 32064 28568 32128
rect 24347 31788 24413 31789
rect 24347 31724 24348 31788
rect 24412 31724 24413 31788
rect 24347 31723 24413 31724
rect 22908 31520 22916 31584
rect 22980 31520 22996 31584
rect 23060 31520 23076 31584
rect 23140 31520 23156 31584
rect 23220 31520 23236 31584
rect 23300 31520 23308 31584
rect 22908 30496 23308 31520
rect 22908 30432 22916 30496
rect 22980 30432 22996 30496
rect 23060 30432 23076 30496
rect 23140 30432 23156 30496
rect 23220 30432 23236 30496
rect 23300 30432 23308 30496
rect 22908 30364 23308 30432
rect 22908 30128 22990 30364
rect 23226 30128 23308 30364
rect 22908 29408 23308 30128
rect 22908 29344 22916 29408
rect 22980 29344 22996 29408
rect 23060 29344 23076 29408
rect 23140 29344 23156 29408
rect 23220 29344 23236 29408
rect 23300 29344 23308 29408
rect 22908 28320 23308 29344
rect 22908 28256 22916 28320
rect 22980 28256 22996 28320
rect 23060 28256 23076 28320
rect 23140 28256 23156 28320
rect 23220 28256 23236 28320
rect 23300 28256 23308 28320
rect 22908 27232 23308 28256
rect 22908 27168 22916 27232
rect 22980 27168 22996 27232
rect 23060 27168 23076 27232
rect 23140 27168 23156 27232
rect 23220 27168 23236 27232
rect 23300 27168 23308 27232
rect 22908 26144 23308 27168
rect 22908 26080 22916 26144
rect 22980 26080 22996 26144
rect 23060 26080 23076 26144
rect 23140 26080 23156 26144
rect 23220 26080 23236 26144
rect 23300 26080 23308 26144
rect 22908 25056 23308 26080
rect 22908 24992 22916 25056
rect 22980 24992 22996 25056
rect 23060 24992 23076 25056
rect 23140 24992 23156 25056
rect 23220 24992 23236 25056
rect 23300 24992 23308 25056
rect 22908 24364 23308 24992
rect 22908 24128 22990 24364
rect 23226 24128 23308 24364
rect 22908 23968 23308 24128
rect 22908 23904 22916 23968
rect 22980 23904 22996 23968
rect 23060 23904 23076 23968
rect 23140 23904 23156 23968
rect 23220 23904 23236 23968
rect 23300 23904 23308 23968
rect 22908 22880 23308 23904
rect 22908 22816 22916 22880
rect 22980 22816 22996 22880
rect 23060 22816 23076 22880
rect 23140 22816 23156 22880
rect 23220 22816 23236 22880
rect 23300 22816 23308 22880
rect 22908 21792 23308 22816
rect 24350 21997 24410 31723
rect 27843 31380 27909 31381
rect 27843 31316 27844 31380
rect 27908 31316 27909 31380
rect 27843 31315 27909 31316
rect 24531 27708 24597 27709
rect 24531 27644 24532 27708
rect 24596 27644 24597 27708
rect 24531 27643 24597 27644
rect 24347 21996 24413 21997
rect 24347 21932 24348 21996
rect 24412 21932 24413 21996
rect 24347 21931 24413 21932
rect 22908 21728 22916 21792
rect 22980 21728 22996 21792
rect 23060 21728 23076 21792
rect 23140 21728 23156 21792
rect 23220 21728 23236 21792
rect 23300 21728 23308 21792
rect 22908 20704 23308 21728
rect 22908 20640 22916 20704
rect 22980 20640 22996 20704
rect 23060 20640 23076 20704
rect 23140 20640 23156 20704
rect 23220 20640 23236 20704
rect 23300 20640 23308 20704
rect 22908 19616 23308 20640
rect 22908 19552 22916 19616
rect 22980 19552 22996 19616
rect 23060 19552 23076 19616
rect 23140 19552 23156 19616
rect 23220 19552 23236 19616
rect 23300 19552 23308 19616
rect 22908 18528 23308 19552
rect 22908 18464 22916 18528
rect 22980 18464 22996 18528
rect 23060 18464 23076 18528
rect 23140 18464 23156 18528
rect 23220 18464 23236 18528
rect 23300 18464 23308 18528
rect 22908 18364 23308 18464
rect 22908 18128 22990 18364
rect 23226 18128 23308 18364
rect 22908 17440 23308 18128
rect 22908 17376 22916 17440
rect 22980 17376 22996 17440
rect 23060 17376 23076 17440
rect 23140 17376 23156 17440
rect 23220 17376 23236 17440
rect 23300 17376 23308 17440
rect 22908 16352 23308 17376
rect 22908 16288 22916 16352
rect 22980 16288 22996 16352
rect 23060 16288 23076 16352
rect 23140 16288 23156 16352
rect 23220 16288 23236 16352
rect 23300 16288 23308 16352
rect 22908 15264 23308 16288
rect 22908 15200 22916 15264
rect 22980 15200 22996 15264
rect 23060 15200 23076 15264
rect 23140 15200 23156 15264
rect 23220 15200 23236 15264
rect 23300 15200 23308 15264
rect 22908 14176 23308 15200
rect 24534 15197 24594 27643
rect 27846 17237 27906 31315
rect 28168 31040 28568 32064
rect 28168 30976 28176 31040
rect 28240 30976 28256 31040
rect 28320 30976 28336 31040
rect 28400 30976 28416 31040
rect 28480 30976 28496 31040
rect 28560 30976 28568 31040
rect 28168 29952 28568 30976
rect 28168 29888 28176 29952
rect 28240 29888 28256 29952
rect 28320 29888 28336 29952
rect 28400 29888 28416 29952
rect 28480 29888 28496 29952
rect 28560 29888 28568 29952
rect 28168 29624 28568 29888
rect 28168 29388 28250 29624
rect 28486 29388 28568 29624
rect 28168 28864 28568 29388
rect 28168 28800 28176 28864
rect 28240 28800 28256 28864
rect 28320 28800 28336 28864
rect 28400 28800 28416 28864
rect 28480 28800 28496 28864
rect 28560 28800 28568 28864
rect 28168 27776 28568 28800
rect 28168 27712 28176 27776
rect 28240 27712 28256 27776
rect 28320 27712 28336 27776
rect 28400 27712 28416 27776
rect 28480 27712 28496 27776
rect 28560 27712 28568 27776
rect 28168 26688 28568 27712
rect 28168 26624 28176 26688
rect 28240 26624 28256 26688
rect 28320 26624 28336 26688
rect 28400 26624 28416 26688
rect 28480 26624 28496 26688
rect 28560 26624 28568 26688
rect 28168 25600 28568 26624
rect 28168 25536 28176 25600
rect 28240 25536 28256 25600
rect 28320 25536 28336 25600
rect 28400 25536 28416 25600
rect 28480 25536 28496 25600
rect 28560 25536 28568 25600
rect 28168 24512 28568 25536
rect 28168 24448 28176 24512
rect 28240 24448 28256 24512
rect 28320 24448 28336 24512
rect 28400 24448 28416 24512
rect 28480 24448 28496 24512
rect 28560 24448 28568 24512
rect 28168 23624 28568 24448
rect 28168 23424 28250 23624
rect 28486 23424 28568 23624
rect 28168 23360 28176 23424
rect 28240 23388 28250 23424
rect 28486 23388 28496 23424
rect 28240 23360 28256 23388
rect 28320 23360 28336 23388
rect 28400 23360 28416 23388
rect 28480 23360 28496 23388
rect 28560 23360 28568 23424
rect 28168 22336 28568 23360
rect 28168 22272 28176 22336
rect 28240 22272 28256 22336
rect 28320 22272 28336 22336
rect 28400 22272 28416 22336
rect 28480 22272 28496 22336
rect 28560 22272 28568 22336
rect 28168 21248 28568 22272
rect 28168 21184 28176 21248
rect 28240 21184 28256 21248
rect 28320 21184 28336 21248
rect 28400 21184 28416 21248
rect 28480 21184 28496 21248
rect 28560 21184 28568 21248
rect 28168 20160 28568 21184
rect 28168 20096 28176 20160
rect 28240 20096 28256 20160
rect 28320 20096 28336 20160
rect 28400 20096 28416 20160
rect 28480 20096 28496 20160
rect 28560 20096 28568 20160
rect 28168 19072 28568 20096
rect 28168 19008 28176 19072
rect 28240 19008 28256 19072
rect 28320 19008 28336 19072
rect 28400 19008 28416 19072
rect 28480 19008 28496 19072
rect 28560 19008 28568 19072
rect 28168 17984 28568 19008
rect 28168 17920 28176 17984
rect 28240 17920 28256 17984
rect 28320 17920 28336 17984
rect 28400 17920 28416 17984
rect 28480 17920 28496 17984
rect 28560 17920 28568 17984
rect 28168 17624 28568 17920
rect 28168 17388 28250 17624
rect 28486 17388 28568 17624
rect 27843 17236 27909 17237
rect 27843 17172 27844 17236
rect 27908 17172 27909 17236
rect 27843 17171 27909 17172
rect 28168 16896 28568 17388
rect 28168 16832 28176 16896
rect 28240 16832 28256 16896
rect 28320 16832 28336 16896
rect 28400 16832 28416 16896
rect 28480 16832 28496 16896
rect 28560 16832 28568 16896
rect 28168 15808 28568 16832
rect 28168 15744 28176 15808
rect 28240 15744 28256 15808
rect 28320 15744 28336 15808
rect 28400 15744 28416 15808
rect 28480 15744 28496 15808
rect 28560 15744 28568 15808
rect 24531 15196 24597 15197
rect 24531 15132 24532 15196
rect 24596 15132 24597 15196
rect 24531 15131 24597 15132
rect 22908 14112 22916 14176
rect 22980 14112 22996 14176
rect 23060 14112 23076 14176
rect 23140 14112 23156 14176
rect 23220 14112 23236 14176
rect 23300 14112 23308 14176
rect 22908 13088 23308 14112
rect 22908 13024 22916 13088
rect 22980 13024 22996 13088
rect 23060 13024 23076 13088
rect 23140 13024 23156 13088
rect 23220 13024 23236 13088
rect 23300 13024 23308 13088
rect 22908 12364 23308 13024
rect 22908 12128 22990 12364
rect 23226 12128 23308 12364
rect 22908 12000 23308 12128
rect 22908 11936 22916 12000
rect 22980 11936 22996 12000
rect 23060 11936 23076 12000
rect 23140 11936 23156 12000
rect 23220 11936 23236 12000
rect 23300 11936 23308 12000
rect 22908 10912 23308 11936
rect 22908 10848 22916 10912
rect 22980 10848 22996 10912
rect 23060 10848 23076 10912
rect 23140 10848 23156 10912
rect 23220 10848 23236 10912
rect 23300 10848 23308 10912
rect 22908 9824 23308 10848
rect 22908 9760 22916 9824
rect 22980 9760 22996 9824
rect 23060 9760 23076 9824
rect 23140 9760 23156 9824
rect 23220 9760 23236 9824
rect 23300 9760 23308 9824
rect 22908 8736 23308 9760
rect 22908 8672 22916 8736
rect 22980 8672 22996 8736
rect 23060 8672 23076 8736
rect 23140 8672 23156 8736
rect 23220 8672 23236 8736
rect 23300 8672 23308 8736
rect 22908 7648 23308 8672
rect 22908 7584 22916 7648
rect 22980 7584 22996 7648
rect 23060 7584 23076 7648
rect 23140 7584 23156 7648
rect 23220 7584 23236 7648
rect 23300 7584 23308 7648
rect 22908 6560 23308 7584
rect 22908 6496 22916 6560
rect 22980 6496 22996 6560
rect 23060 6496 23076 6560
rect 23140 6496 23156 6560
rect 23220 6496 23236 6560
rect 23300 6496 23308 6560
rect 22908 6364 23308 6496
rect 22908 6128 22990 6364
rect 23226 6128 23308 6364
rect 22908 5472 23308 6128
rect 22908 5408 22916 5472
rect 22980 5408 22996 5472
rect 23060 5408 23076 5472
rect 23140 5408 23156 5472
rect 23220 5408 23236 5472
rect 23300 5408 23308 5472
rect 22908 4384 23308 5408
rect 22908 4320 22916 4384
rect 22980 4320 22996 4384
rect 23060 4320 23076 4384
rect 23140 4320 23156 4384
rect 23220 4320 23236 4384
rect 23300 4320 23308 4384
rect 22908 3296 23308 4320
rect 22908 3232 22916 3296
rect 22980 3232 22996 3296
rect 23060 3232 23076 3296
rect 23140 3232 23156 3296
rect 23220 3232 23236 3296
rect 23300 3232 23308 3296
rect 22908 2208 23308 3232
rect 22908 2144 22916 2208
rect 22980 2144 22996 2208
rect 23060 2144 23076 2208
rect 23140 2144 23156 2208
rect 23220 2144 23236 2208
rect 23300 2144 23308 2208
rect 22908 2128 23308 2144
rect 28168 14720 28568 15744
rect 28168 14656 28176 14720
rect 28240 14656 28256 14720
rect 28320 14656 28336 14720
rect 28400 14656 28416 14720
rect 28480 14656 28496 14720
rect 28560 14656 28568 14720
rect 28168 13632 28568 14656
rect 28168 13568 28176 13632
rect 28240 13568 28256 13632
rect 28320 13568 28336 13632
rect 28400 13568 28416 13632
rect 28480 13568 28496 13632
rect 28560 13568 28568 13632
rect 28168 12544 28568 13568
rect 28168 12480 28176 12544
rect 28240 12480 28256 12544
rect 28320 12480 28336 12544
rect 28400 12480 28416 12544
rect 28480 12480 28496 12544
rect 28560 12480 28568 12544
rect 28168 11624 28568 12480
rect 28168 11456 28250 11624
rect 28486 11456 28568 11624
rect 28168 11392 28176 11456
rect 28240 11392 28250 11456
rect 28486 11392 28496 11456
rect 28560 11392 28568 11456
rect 28168 11388 28250 11392
rect 28486 11388 28568 11392
rect 28168 10368 28568 11388
rect 28168 10304 28176 10368
rect 28240 10304 28256 10368
rect 28320 10304 28336 10368
rect 28400 10304 28416 10368
rect 28480 10304 28496 10368
rect 28560 10304 28568 10368
rect 28168 9280 28568 10304
rect 28168 9216 28176 9280
rect 28240 9216 28256 9280
rect 28320 9216 28336 9280
rect 28400 9216 28416 9280
rect 28480 9216 28496 9280
rect 28560 9216 28568 9280
rect 28168 8192 28568 9216
rect 28168 8128 28176 8192
rect 28240 8128 28256 8192
rect 28320 8128 28336 8192
rect 28400 8128 28416 8192
rect 28480 8128 28496 8192
rect 28560 8128 28568 8192
rect 28168 7104 28568 8128
rect 28168 7040 28176 7104
rect 28240 7040 28256 7104
rect 28320 7040 28336 7104
rect 28400 7040 28416 7104
rect 28480 7040 28496 7104
rect 28560 7040 28568 7104
rect 28168 6016 28568 7040
rect 28168 5952 28176 6016
rect 28240 5952 28256 6016
rect 28320 5952 28336 6016
rect 28400 5952 28416 6016
rect 28480 5952 28496 6016
rect 28560 5952 28568 6016
rect 28168 5624 28568 5952
rect 28168 5388 28250 5624
rect 28486 5388 28568 5624
rect 28168 4928 28568 5388
rect 28168 4864 28176 4928
rect 28240 4864 28256 4928
rect 28320 4864 28336 4928
rect 28400 4864 28416 4928
rect 28480 4864 28496 4928
rect 28560 4864 28568 4928
rect 28168 3840 28568 4864
rect 28168 3776 28176 3840
rect 28240 3776 28256 3840
rect 28320 3776 28336 3840
rect 28400 3776 28416 3840
rect 28480 3776 28496 3840
rect 28560 3776 28568 3840
rect 28168 2752 28568 3776
rect 28168 2688 28176 2752
rect 28240 2688 28256 2752
rect 28320 2688 28336 2752
rect 28400 2688 28416 2752
rect 28480 2688 28496 2752
rect 28560 2688 28568 2752
rect 28168 2128 28568 2688
rect 28908 31584 29308 32144
rect 28908 31520 28916 31584
rect 28980 31520 28996 31584
rect 29060 31520 29076 31584
rect 29140 31520 29156 31584
rect 29220 31520 29236 31584
rect 29300 31520 29308 31584
rect 28908 30496 29308 31520
rect 28908 30432 28916 30496
rect 28980 30432 28996 30496
rect 29060 30432 29076 30496
rect 29140 30432 29156 30496
rect 29220 30432 29236 30496
rect 29300 30432 29308 30496
rect 28908 30364 29308 30432
rect 28908 30128 28990 30364
rect 29226 30128 29308 30364
rect 28908 29408 29308 30128
rect 28908 29344 28916 29408
rect 28980 29344 28996 29408
rect 29060 29344 29076 29408
rect 29140 29344 29156 29408
rect 29220 29344 29236 29408
rect 29300 29344 29308 29408
rect 28908 28320 29308 29344
rect 28908 28256 28916 28320
rect 28980 28256 28996 28320
rect 29060 28256 29076 28320
rect 29140 28256 29156 28320
rect 29220 28256 29236 28320
rect 29300 28256 29308 28320
rect 28908 27232 29308 28256
rect 28908 27168 28916 27232
rect 28980 27168 28996 27232
rect 29060 27168 29076 27232
rect 29140 27168 29156 27232
rect 29220 27168 29236 27232
rect 29300 27168 29308 27232
rect 28908 26144 29308 27168
rect 28908 26080 28916 26144
rect 28980 26080 28996 26144
rect 29060 26080 29076 26144
rect 29140 26080 29156 26144
rect 29220 26080 29236 26144
rect 29300 26080 29308 26144
rect 28908 25056 29308 26080
rect 28908 24992 28916 25056
rect 28980 24992 28996 25056
rect 29060 24992 29076 25056
rect 29140 24992 29156 25056
rect 29220 24992 29236 25056
rect 29300 24992 29308 25056
rect 28908 24364 29308 24992
rect 28908 24128 28990 24364
rect 29226 24128 29308 24364
rect 28908 23968 29308 24128
rect 28908 23904 28916 23968
rect 28980 23904 28996 23968
rect 29060 23904 29076 23968
rect 29140 23904 29156 23968
rect 29220 23904 29236 23968
rect 29300 23904 29308 23968
rect 28908 22880 29308 23904
rect 28908 22816 28916 22880
rect 28980 22816 28996 22880
rect 29060 22816 29076 22880
rect 29140 22816 29156 22880
rect 29220 22816 29236 22880
rect 29300 22816 29308 22880
rect 28908 21792 29308 22816
rect 28908 21728 28916 21792
rect 28980 21728 28996 21792
rect 29060 21728 29076 21792
rect 29140 21728 29156 21792
rect 29220 21728 29236 21792
rect 29300 21728 29308 21792
rect 28908 20704 29308 21728
rect 28908 20640 28916 20704
rect 28980 20640 28996 20704
rect 29060 20640 29076 20704
rect 29140 20640 29156 20704
rect 29220 20640 29236 20704
rect 29300 20640 29308 20704
rect 28908 19616 29308 20640
rect 28908 19552 28916 19616
rect 28980 19552 28996 19616
rect 29060 19552 29076 19616
rect 29140 19552 29156 19616
rect 29220 19552 29236 19616
rect 29300 19552 29308 19616
rect 28908 18528 29308 19552
rect 28908 18464 28916 18528
rect 28980 18464 28996 18528
rect 29060 18464 29076 18528
rect 29140 18464 29156 18528
rect 29220 18464 29236 18528
rect 29300 18464 29308 18528
rect 28908 18364 29308 18464
rect 28908 18128 28990 18364
rect 29226 18128 29308 18364
rect 28908 17440 29308 18128
rect 28908 17376 28916 17440
rect 28980 17376 28996 17440
rect 29060 17376 29076 17440
rect 29140 17376 29156 17440
rect 29220 17376 29236 17440
rect 29300 17376 29308 17440
rect 28908 16352 29308 17376
rect 28908 16288 28916 16352
rect 28980 16288 28996 16352
rect 29060 16288 29076 16352
rect 29140 16288 29156 16352
rect 29220 16288 29236 16352
rect 29300 16288 29308 16352
rect 28908 15264 29308 16288
rect 28908 15200 28916 15264
rect 28980 15200 28996 15264
rect 29060 15200 29076 15264
rect 29140 15200 29156 15264
rect 29220 15200 29236 15264
rect 29300 15200 29308 15264
rect 28908 14176 29308 15200
rect 28908 14112 28916 14176
rect 28980 14112 28996 14176
rect 29060 14112 29076 14176
rect 29140 14112 29156 14176
rect 29220 14112 29236 14176
rect 29300 14112 29308 14176
rect 28908 13088 29308 14112
rect 28908 13024 28916 13088
rect 28980 13024 28996 13088
rect 29060 13024 29076 13088
rect 29140 13024 29156 13088
rect 29220 13024 29236 13088
rect 29300 13024 29308 13088
rect 28908 12364 29308 13024
rect 28908 12128 28990 12364
rect 29226 12128 29308 12364
rect 28908 12000 29308 12128
rect 28908 11936 28916 12000
rect 28980 11936 28996 12000
rect 29060 11936 29076 12000
rect 29140 11936 29156 12000
rect 29220 11936 29236 12000
rect 29300 11936 29308 12000
rect 28908 10912 29308 11936
rect 28908 10848 28916 10912
rect 28980 10848 28996 10912
rect 29060 10848 29076 10912
rect 29140 10848 29156 10912
rect 29220 10848 29236 10912
rect 29300 10848 29308 10912
rect 28908 9824 29308 10848
rect 28908 9760 28916 9824
rect 28980 9760 28996 9824
rect 29060 9760 29076 9824
rect 29140 9760 29156 9824
rect 29220 9760 29236 9824
rect 29300 9760 29308 9824
rect 28908 8736 29308 9760
rect 28908 8672 28916 8736
rect 28980 8672 28996 8736
rect 29060 8672 29076 8736
rect 29140 8672 29156 8736
rect 29220 8672 29236 8736
rect 29300 8672 29308 8736
rect 28908 7648 29308 8672
rect 28908 7584 28916 7648
rect 28980 7584 28996 7648
rect 29060 7584 29076 7648
rect 29140 7584 29156 7648
rect 29220 7584 29236 7648
rect 29300 7584 29308 7648
rect 28908 6560 29308 7584
rect 28908 6496 28916 6560
rect 28980 6496 28996 6560
rect 29060 6496 29076 6560
rect 29140 6496 29156 6560
rect 29220 6496 29236 6560
rect 29300 6496 29308 6560
rect 28908 6364 29308 6496
rect 28908 6128 28990 6364
rect 29226 6128 29308 6364
rect 28908 5472 29308 6128
rect 28908 5408 28916 5472
rect 28980 5408 28996 5472
rect 29060 5408 29076 5472
rect 29140 5408 29156 5472
rect 29220 5408 29236 5472
rect 29300 5408 29308 5472
rect 28908 4384 29308 5408
rect 28908 4320 28916 4384
rect 28980 4320 28996 4384
rect 29060 4320 29076 4384
rect 29140 4320 29156 4384
rect 29220 4320 29236 4384
rect 29300 4320 29308 4384
rect 28908 3296 29308 4320
rect 28908 3232 28916 3296
rect 28980 3232 28996 3296
rect 29060 3232 29076 3296
rect 29140 3232 29156 3296
rect 29220 3232 29236 3296
rect 29300 3232 29308 3296
rect 28908 2208 29308 3232
rect 28908 2144 28916 2208
rect 28980 2144 28996 2208
rect 29060 2144 29076 2208
rect 29140 2144 29156 2208
rect 29220 2144 29236 2208
rect 29300 2144 29308 2208
rect 28908 2128 29308 2144
<< via4 >>
rect 4250 29388 4486 29624
rect 4250 23424 4486 23624
rect 4250 23388 4256 23424
rect 4256 23388 4320 23424
rect 4320 23388 4336 23424
rect 4336 23388 4400 23424
rect 4400 23388 4416 23424
rect 4416 23388 4480 23424
rect 4480 23388 4486 23424
rect 4250 17388 4486 17624
rect 4250 11456 4486 11624
rect 4250 11392 4256 11456
rect 4256 11392 4320 11456
rect 4320 11392 4336 11456
rect 4336 11392 4400 11456
rect 4400 11392 4416 11456
rect 4416 11392 4480 11456
rect 4480 11392 4486 11456
rect 4250 11388 4486 11392
rect 4250 5388 4486 5624
rect 4990 30128 5226 30364
rect 4990 24128 5226 24364
rect 4990 18128 5226 18364
rect 4990 12128 5226 12364
rect 4990 6128 5226 6364
rect 10250 29388 10486 29624
rect 10250 23424 10486 23624
rect 10250 23388 10256 23424
rect 10256 23388 10320 23424
rect 10320 23388 10336 23424
rect 10336 23388 10400 23424
rect 10400 23388 10416 23424
rect 10416 23388 10480 23424
rect 10480 23388 10486 23424
rect 10250 17388 10486 17624
rect 10250 11456 10486 11624
rect 10250 11392 10256 11456
rect 10256 11392 10320 11456
rect 10320 11392 10336 11456
rect 10336 11392 10400 11456
rect 10400 11392 10416 11456
rect 10416 11392 10480 11456
rect 10480 11392 10486 11456
rect 10250 11388 10486 11392
rect 10250 5388 10486 5624
rect 10990 30128 11226 30364
rect 10990 24128 11226 24364
rect 16250 29388 16486 29624
rect 10990 18128 11226 18364
rect 16250 23424 16486 23624
rect 16250 23388 16256 23424
rect 16256 23388 16320 23424
rect 16320 23388 16336 23424
rect 16336 23388 16400 23424
rect 16400 23388 16416 23424
rect 16416 23388 16480 23424
rect 16480 23388 16486 23424
rect 16250 17388 16486 17624
rect 10990 12128 11226 12364
rect 16250 11456 16486 11624
rect 16250 11392 16256 11456
rect 16256 11392 16320 11456
rect 16320 11392 16336 11456
rect 16336 11392 16400 11456
rect 16400 11392 16416 11456
rect 16416 11392 16480 11456
rect 16480 11392 16486 11456
rect 16250 11388 16486 11392
rect 10990 6128 11226 6364
rect 16250 5388 16486 5624
rect 16990 30128 17226 30364
rect 22250 29388 22486 29624
rect 16990 24128 17226 24364
rect 16990 18128 17226 18364
rect 16990 12128 17226 12364
rect 22250 23424 22486 23624
rect 22250 23388 22256 23424
rect 22256 23388 22320 23424
rect 22320 23388 22336 23424
rect 22336 23388 22400 23424
rect 22400 23388 22416 23424
rect 22416 23388 22480 23424
rect 22480 23388 22486 23424
rect 22250 17388 22486 17624
rect 22250 11456 22486 11624
rect 22250 11392 22256 11456
rect 22256 11392 22320 11456
rect 22320 11392 22336 11456
rect 22336 11392 22400 11456
rect 22400 11392 22416 11456
rect 22416 11392 22480 11456
rect 22480 11392 22486 11456
rect 22250 11388 22486 11392
rect 16990 6128 17226 6364
rect 22250 5388 22486 5624
rect 22990 30128 23226 30364
rect 22990 24128 23226 24364
rect 22990 18128 23226 18364
rect 28250 29388 28486 29624
rect 28250 23424 28486 23624
rect 28250 23388 28256 23424
rect 28256 23388 28320 23424
rect 28320 23388 28336 23424
rect 28336 23388 28400 23424
rect 28400 23388 28416 23424
rect 28416 23388 28480 23424
rect 28480 23388 28486 23424
rect 28250 17388 28486 17624
rect 22990 12128 23226 12364
rect 22990 6128 23226 6364
rect 28250 11456 28486 11624
rect 28250 11392 28256 11456
rect 28256 11392 28320 11456
rect 28320 11392 28336 11456
rect 28336 11392 28400 11456
rect 28400 11392 28416 11456
rect 28416 11392 28480 11456
rect 28480 11392 28486 11456
rect 28250 11388 28486 11392
rect 28250 5388 28486 5624
rect 28990 30128 29226 30364
rect 28990 24128 29226 24364
rect 28990 18128 29226 18364
rect 28990 12128 29226 12364
rect 28990 6128 29226 6364
<< metal5 >>
rect 1056 30364 31328 30446
rect 1056 30128 4990 30364
rect 5226 30128 10990 30364
rect 11226 30128 16990 30364
rect 17226 30128 22990 30364
rect 23226 30128 28990 30364
rect 29226 30128 31328 30364
rect 1056 30046 31328 30128
rect 1056 29624 31328 29706
rect 1056 29388 4250 29624
rect 4486 29388 10250 29624
rect 10486 29388 16250 29624
rect 16486 29388 22250 29624
rect 22486 29388 28250 29624
rect 28486 29388 31328 29624
rect 1056 29306 31328 29388
rect 1056 24364 31328 24446
rect 1056 24128 4990 24364
rect 5226 24128 10990 24364
rect 11226 24128 16990 24364
rect 17226 24128 22990 24364
rect 23226 24128 28990 24364
rect 29226 24128 31328 24364
rect 1056 24046 31328 24128
rect 1056 23624 31328 23706
rect 1056 23388 4250 23624
rect 4486 23388 10250 23624
rect 10486 23388 16250 23624
rect 16486 23388 22250 23624
rect 22486 23388 28250 23624
rect 28486 23388 31328 23624
rect 1056 23306 31328 23388
rect 1056 18364 31328 18446
rect 1056 18128 4990 18364
rect 5226 18128 10990 18364
rect 11226 18128 16990 18364
rect 17226 18128 22990 18364
rect 23226 18128 28990 18364
rect 29226 18128 31328 18364
rect 1056 18046 31328 18128
rect 1056 17624 31328 17706
rect 1056 17388 4250 17624
rect 4486 17388 10250 17624
rect 10486 17388 16250 17624
rect 16486 17388 22250 17624
rect 22486 17388 28250 17624
rect 28486 17388 31328 17624
rect 1056 17306 31328 17388
rect 1056 12364 31328 12446
rect 1056 12128 4990 12364
rect 5226 12128 10990 12364
rect 11226 12128 16990 12364
rect 17226 12128 22990 12364
rect 23226 12128 28990 12364
rect 29226 12128 31328 12364
rect 1056 12046 31328 12128
rect 1056 11624 31328 11706
rect 1056 11388 4250 11624
rect 4486 11388 10250 11624
rect 10486 11388 16250 11624
rect 16486 11388 22250 11624
rect 22486 11388 28250 11624
rect 28486 11388 31328 11624
rect 1056 11306 31328 11388
rect 1056 6364 31328 6446
rect 1056 6128 4990 6364
rect 5226 6128 10990 6364
rect 11226 6128 16990 6364
rect 17226 6128 22990 6364
rect 23226 6128 28990 6364
rect 29226 6128 31328 6364
rect 1056 6046 31328 6128
rect 1056 5624 31328 5706
rect 1056 5388 4250 5624
rect 4486 5388 10250 5624
rect 10486 5388 16250 5624
rect 16486 5388 22250 5624
rect 22486 5388 28250 5624
rect 28486 5388 31328 5624
rect 1056 5306 31328 5388
use sky130_fd_sc_hd__or4_4  _0480_
timestamp 0
transform 1 0 24656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0481_
timestamp 0
transform 1 0 18400 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0482_
timestamp 0
transform -1 0 25024 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor4_1  _0483_
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0484_
timestamp 0
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _0485_
timestamp 0
transform -1 0 24012 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0486_
timestamp 0
transform -1 0 24748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0487_
timestamp 0
transform -1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0488_
timestamp 0
transform -1 0 22080 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0489_
timestamp 0
transform -1 0 22540 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0490_
timestamp 0
transform -1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0491_
timestamp 0
transform 1 0 24288 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0492_
timestamp 0
transform 1 0 25024 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0493_
timestamp 0
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0494_
timestamp 0
transform -1 0 21344 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0495_
timestamp 0
transform -1 0 14904 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0496_
timestamp 0
transform 1 0 22908 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0497_
timestamp 0
transform 1 0 23736 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0498_
timestamp 0
transform -1 0 23184 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0499_
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_4  _0500_
timestamp 0
transform 1 0 20424 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0501_
timestamp 0
transform 1 0 21252 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0502_
timestamp 0
transform -1 0 21712 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0503_
timestamp 0
transform -1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0504_
timestamp 0
transform -1 0 20240 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_4  _0505_
timestamp 0
transform 1 0 20240 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0506_
timestamp 0
transform 1 0 18492 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0507_
timestamp 0
transform 1 0 20700 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_1  _0508_
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0509_
timestamp 0
transform 1 0 23368 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0510_
timestamp 0
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0511_
timestamp 0
transform -1 0 24288 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0512_
timestamp 0
transform 1 0 20516 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and4bb_4  _0513_
timestamp 0
transform 1 0 20516 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0514_
timestamp 0
transform 1 0 19688 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0515_
timestamp 0
transform 1 0 23092 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4b_2  _0516_
timestamp 0
transform -1 0 24196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _0517_
timestamp 0
transform 1 0 23736 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_2  _0518_
timestamp 0
transform -1 0 23092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__and4b_1  _0519_
timestamp 0
transform 1 0 21712 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0520_
timestamp 0
transform -1 0 22356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0521_
timestamp 0
transform 1 0 21804 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0522_
timestamp 0
transform 1 0 22540 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0523_
timestamp 0
transform 1 0 24380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0524_
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0525_
timestamp 0
transform 1 0 19688 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0526_
timestamp 0
transform -1 0 18400 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0527_
timestamp 0
transform -1 0 20424 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0528_
timestamp 0
transform -1 0 26956 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0529_
timestamp 0
transform 1 0 26680 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0530_
timestamp 0
transform 1 0 22908 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0531_
timestamp 0
transform 1 0 23552 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0532_
timestamp 0
transform 1 0 18124 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0533_
timestamp 0
transform 1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0534_
timestamp 0
transform -1 0 24656 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0535_
timestamp 0
transform 1 0 19412 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0536_
timestamp 0
transform 1 0 24104 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0537_
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0538_
timestamp 0
transform 1 0 23552 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0539_
timestamp 0
transform 1 0 24380 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0540_
timestamp 0
transform 1 0 25484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 0
transform 1 0 26128 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0542_
timestamp 0
transform -1 0 11776 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0543_
timestamp 0
transform 1 0 10488 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0544_
timestamp 0
transform 1 0 4416 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0545_
timestamp 0
transform 1 0 7912 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0546_
timestamp 0
transform 1 0 10120 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0547_
timestamp 0
transform -1 0 12972 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0548_
timestamp 0
transform 1 0 12420 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0549_
timestamp 0
transform 1 0 6992 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0550_
timestamp 0
transform 1 0 10672 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0551_
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0552_
timestamp 0
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0553_
timestamp 0
transform -1 0 12512 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0554_
timestamp 0
transform 1 0 22172 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 0
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0556_
timestamp 0
transform 1 0 17756 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0557_
timestamp 0
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0558_
timestamp 0
transform 1 0 22816 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0559_
timestamp 0
transform 1 0 19504 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0560_
timestamp 0
transform 1 0 23552 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0561_
timestamp 0
transform 1 0 22816 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0562_
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0563_
timestamp 0
transform 1 0 25116 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0564_
timestamp 0
transform -1 0 27508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 0
transform 1 0 26036 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0566_
timestamp 0
transform 1 0 10672 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0567_
timestamp 0
transform 1 0 10580 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0568_
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0569_
timestamp 0
transform 1 0 5796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0570_
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0571_
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0572_
timestamp 0
transform 1 0 13340 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0573_
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0574_
timestamp 0
transform -1 0 12052 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0575_
timestamp 0
transform 1 0 11316 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0576_
timestamp 0
transform -1 0 15456 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0577_
timestamp 0
transform -1 0 12696 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0578_
timestamp 0
transform 1 0 10672 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0579_
timestamp 0
transform 1 0 11316 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0580_
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0581_
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0582_
timestamp 0
transform 1 0 10488 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp 0
transform 1 0 11592 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0584_
timestamp 0
transform 1 0 12328 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0585_
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0586_
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0587_
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0588_
timestamp 0
transform -1 0 15548 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 0
transform 1 0 11684 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0590_
timestamp 0
transform 1 0 10948 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0591_
timestamp 0
transform 1 0 11592 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp 0
transform 1 0 4784 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0593_
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0594_
timestamp 0
transform 1 0 10488 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0595_
timestamp 0
transform -1 0 14996 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0596_
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp 0
transform 1 0 7176 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0598_
timestamp 0
transform 1 0 11592 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0599_
timestamp 0
transform 1 0 12236 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0600_
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0601_
timestamp 0
transform 1 0 12696 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0602_
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0603_
timestamp 0
transform 1 0 15364 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp 0
transform 1 0 4968 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0605_
timestamp 0
transform 1 0 7912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 0
transform 1 0 12052 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0607_
timestamp 0
transform 1 0 14904 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0608_
timestamp 0
transform 1 0 16376 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0609_
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0610_
timestamp 0
transform 1 0 15548 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0611_
timestamp 0
transform 1 0 16100 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0612_
timestamp 0
transform -1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0613_
timestamp 0
transform 1 0 17020 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0614_
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0615_
timestamp 0
transform -1 0 18032 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0616_
timestamp 0
transform 1 0 18032 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0617_
timestamp 0
transform 1 0 17480 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0618_
timestamp 0
transform -1 0 23552 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0619_
timestamp 0
transform -1 0 23000 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0620_
timestamp 0
transform 1 0 18400 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0621_
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0622_
timestamp 0
transform -1 0 20056 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0623_
timestamp 0
transform 1 0 20792 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0624_
timestamp 0
transform -1 0 19504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0625_
timestamp 0
transform 1 0 20056 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 0
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 0
transform -1 0 18768 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0628_
timestamp 0
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0629_
timestamp 0
transform -1 0 19044 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0630_
timestamp 0
transform -1 0 24012 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0631_
timestamp 0
transform -1 0 25392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 0
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0633_
timestamp 0
transform -1 0 25024 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0634_
timestamp 0
transform 1 0 22724 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0635_
timestamp 0
transform 1 0 24104 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0636_
timestamp 0
transform -1 0 25300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0637_
timestamp 0
transform -1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0638_
timestamp 0
transform -1 0 23736 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0639_
timestamp 0
transform -1 0 24472 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0640_
timestamp 0
transform -1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0641_
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 0
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0643_
timestamp 0
transform 1 0 20884 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0644_
timestamp 0
transform -1 0 21252 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0645_
timestamp 0
transform -1 0 19596 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _0646_
timestamp 0
transform 1 0 7912 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 0
transform -1 0 22080 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0648_
timestamp 0
transform 1 0 20516 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0649_
timestamp 0
transform 1 0 14812 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0650_
timestamp 0
transform -1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0651_
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0652_
timestamp 0
transform 1 0 12328 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0653_
timestamp 0
transform -1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0654_
timestamp 0
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0655_
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0656_
timestamp 0
transform -1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0657_
timestamp 0
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 0
transform -1 0 11224 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 0
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0660_
timestamp 0
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0661_
timestamp 0
transform 1 0 24196 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0662_
timestamp 0
transform -1 0 24196 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0663_
timestamp 0
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0664_
timestamp 0
transform 1 0 10672 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0665_
timestamp 0
transform 1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0666_
timestamp 0
transform -1 0 26864 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0667_
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0668_
timestamp 0
transform -1 0 23828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0669_
timestamp 0
transform 1 0 26128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0670_
timestamp 0
transform -1 0 25300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0671_
timestamp 0
transform 1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0672_
timestamp 0
transform -1 0 27784 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 0
transform -1 0 27232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 0
transform 1 0 27048 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 0
transform -1 0 26772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 0
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0678_
timestamp 0
transform -1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 0
transform -1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0680_
timestamp 0
transform -1 0 15088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 0
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 0
transform 1 0 27140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0683_
timestamp 0
transform -1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 0
transform -1 0 29532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 0
transform -1 0 28704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0686_
timestamp 0
transform -1 0 18584 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  _0687_
timestamp 0
transform -1 0 17848 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__a21o_1  _0688_
timestamp 0
transform 1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0689_
timestamp 0
transform -1 0 17572 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0690_
timestamp 0
transform 1 0 16008 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0691_
timestamp 0
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0693_
timestamp 0
transform -1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0694_
timestamp 0
transform 1 0 13064 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0695_
timestamp 0
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0696_
timestamp 0
transform -1 0 13892 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0697_
timestamp 0
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0698_
timestamp 0
transform 1 0 25852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0699_
timestamp 0
transform -1 0 25392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0700_
timestamp 0
transform 1 0 12788 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0701_
timestamp 0
transform -1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0702_
timestamp 0
transform -1 0 26864 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0703_
timestamp 0
transform -1 0 27232 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 0
transform 1 0 26036 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0705_
timestamp 0
transform -1 0 26036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0706_
timestamp 0
transform -1 0 19136 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0708_
timestamp 0
transform -1 0 16744 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0709_
timestamp 0
transform 1 0 14536 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0710_
timestamp 0
transform -1 0 13984 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0711_
timestamp 0
transform 1 0 13432 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0712_
timestamp 0
transform -1 0 11408 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0713_
timestamp 0
transform 1 0 10488 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0714_
timestamp 0
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0715_
timestamp 0
transform 1 0 8832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0716_
timestamp 0
transform -1 0 8832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0717_
timestamp 0
transform -1 0 24196 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0718_
timestamp 0
transform 1 0 23644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 0
transform 1 0 10212 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0720_
timestamp 0
transform -1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 0
transform 1 0 25300 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0722_
timestamp 0
transform -1 0 23552 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 0
transform -1 0 26128 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0724_
timestamp 0
transform 1 0 26128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0725_
timestamp 0
transform -1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0726_
timestamp 0
transform 1 0 15456 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0727_
timestamp 0
transform -1 0 17388 0 1 17408
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0728_
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0729_
timestamp 0
transform -1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0730_
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0731_
timestamp 0
transform -1 0 5704 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 0
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0733_
timestamp 0
transform -1 0 5428 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0735_
timestamp 0
transform 1 0 5336 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0737_
timestamp 0
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0739_
timestamp 0
transform -1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 0
transform -1 0 19136 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0741_
timestamp 0
transform 1 0 20976 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 0
transform 1 0 19412 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0743_
timestamp 0
transform -1 0 19136 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 0
transform 1 0 15732 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0745_
timestamp 0
transform 1 0 15916 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 0
transform 1 0 6992 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0747_
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 0
transform 1 0 6256 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0749_
timestamp 0
transform 1 0 5336 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0751_
timestamp 0
transform 1 0 5520 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 0
transform 1 0 6532 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0753_
timestamp 0
transform 1 0 5428 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 0
transform -1 0 22080 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0755_
timestamp 0
transform 1 0 22540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 0
transform 1 0 6164 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0757_
timestamp 0
transform -1 0 6164 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 0
transform 1 0 20424 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0759_
timestamp 0
transform -1 0 20056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 0
transform 1 0 21344 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0761_
timestamp 0
transform 1 0 21160 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0762_
timestamp 0
transform 1 0 15272 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0763_
timestamp 0
transform 1 0 15732 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0765_
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 0
transform 1 0 6532 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0767_
timestamp 0
transform -1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0769_
timestamp 0
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 0
transform 1 0 6532 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0771_
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0773_
timestamp 0
transform -1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0775_
timestamp 0
transform 1 0 5888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 0
transform -1 0 19964 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0777_
timestamp 0
transform 1 0 20700 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 0
transform -1 0 20148 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0779_
timestamp 0
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 0
transform -1 0 16376 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0781_
timestamp 0
transform 1 0 15364 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 0
transform -1 0 16560 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0783_
timestamp 0
transform 1 0 16928 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 0
transform 1 0 12972 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0785_
timestamp 0
transform -1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 0
transform 1 0 13340 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0787_
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 0
transform 1 0 13064 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0789_
timestamp 0
transform -1 0 12880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 0
transform 1 0 24196 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0791_
timestamp 0
transform -1 0 24288 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 0
transform 1 0 12696 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0793_
timestamp 0
transform -1 0 12236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 0
transform -1 0 25576 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0795_
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 0
transform -1 0 26036 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0797_
timestamp 0
transform 1 0 26496 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 0
transform 1 0 15732 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _0799_
timestamp 0
transform 1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0801_
timestamp 0
transform 1 0 12696 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 0
transform 1 0 10028 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0803_
timestamp 0
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 0
transform 1 0 9660 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0805_
timestamp 0
transform 1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 0
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0807_
timestamp 0
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0809_
timestamp 0
transform -1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 0
transform 1 0 10212 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0811_
timestamp 0
transform 1 0 9108 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 0
transform 1 0 22080 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0813_
timestamp 0
transform -1 0 21712 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 0
transform -1 0 24012 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0815_
timestamp 0
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0816_
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 0
transform -1 0 19688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0818_
timestamp 0
transform 1 0 18676 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0819_
timestamp 0
transform 1 0 19320 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0821_
timestamp 0
transform 1 0 10488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0822_
timestamp 0
transform 1 0 9476 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0823_
timestamp 0
transform 1 0 8372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0824_
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0825_
timestamp 0
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0826_
timestamp 0
transform 1 0 9292 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0827_
timestamp 0
transform -1 0 8832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0828_
timestamp 0
transform 1 0 23460 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0829_
timestamp 0
transform -1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0831_
timestamp 0
transform 1 0 8280 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0832_
timestamp 0
transform -1 0 25484 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0833_
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0834_
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0835_
timestamp 0
transform -1 0 24288 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0836_
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0837_
timestamp 0
transform -1 0 18032 0 1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0838_
timestamp 0
transform 1 0 14996 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0839_
timestamp 0
transform -1 0 14904 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0840_
timestamp 0
transform 1 0 13892 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0841_
timestamp 0
transform -1 0 13892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 0
transform 1 0 13156 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0843_
timestamp 0
transform 1 0 12512 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 0
transform 1 0 12512 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0845_
timestamp 0
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0847_
timestamp 0
transform -1 0 17480 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 0
transform 1 0 13064 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0849_
timestamp 0
transform -1 0 13064 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 0
transform 1 0 17940 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 0
transform 1 0 17664 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 0
transform 1 0 18308 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0853_
timestamp 0
transform -1 0 17664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 0
transform -1 0 16284 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0855_
timestamp 0
transform 1 0 15272 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 0
transform 1 0 13984 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0857_
timestamp 0
transform -1 0 13984 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 0
transform -1 0 15824 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 0
transform 1 0 16192 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 0
transform 1 0 9384 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 0
transform -1 0 9568 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 0
transform 1 0 9568 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0863_
timestamp 0
transform -1 0 9568 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 0
transform 1 0 18400 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0865_
timestamp 0
transform -1 0 17020 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0866_
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0867_
timestamp 0
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0868_
timestamp 0
transform 1 0 17572 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0869_
timestamp 0
transform -1 0 17296 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 0
transform 1 0 17480 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0871_
timestamp 0
transform 1 0 17204 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0872_
timestamp 0
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0873_
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0874_
timestamp 0
transform 1 0 3404 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 0
transform -1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 0
transform 1 0 4784 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0877_
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0878_
timestamp 0
transform 1 0 3864 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0879_
timestamp 0
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0880_
timestamp 0
transform 1 0 2576 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 0
transform -1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 0
transform 1 0 16192 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0883_
timestamp 0
transform -1 0 14720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0885_
timestamp 0
transform 1 0 2576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 0
transform 1 0 16652 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 0
transform -1 0 16560 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 0
transform 1 0 16744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0889_
timestamp 0
transform -1 0 16192 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 0
transform 1 0 15640 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0891_
timestamp 0
transform -1 0 17940 0 -1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 0
transform 1 0 2576 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 0
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0894_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 0
transform 1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 0
transform 1 0 2576 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 0
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 0
transform 1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0900_
timestamp 0
transform 1 0 15272 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 0
transform 1 0 14996 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0904_
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 0
transform 1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 0
transform 1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0907_
timestamp 0
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0908_
timestamp 0
transform -1 0 18400 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0909_
timestamp 0
transform 1 0 16652 0 1 20672
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 0
transform -1 0 11224 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0912_
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0913_
timestamp 0
transform 1 0 7820 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 0
transform 1 0 7820 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 0
transform 1 0 10120 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 0
transform -1 0 21620 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 0
transform 1 0 8096 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 0
transform -1 0 24288 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 0
transform -1 0 24104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 0
transform 1 0 23092 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 0
transform 1 0 22908 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 0
transform -1 0 17112 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0927_
timestamp 0
transform -1 0 18400 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 0
transform -1 0 5704 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0930_
timestamp 0
transform 1 0 4600 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 0
transform 1 0 4232 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0932_
timestamp 0
transform 1 0 5244 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 0
transform 1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0934_
timestamp 0
transform 1 0 4232 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 0
transform 1 0 3956 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0936_
timestamp 0
transform 1 0 20792 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 0
transform 1 0 20792 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0938_
timestamp 0
transform 1 0 5336 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 0
transform 1 0 4232 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0940_
timestamp 0
transform 1 0 20608 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 0
transform 1 0 20516 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0942_
timestamp 0
transform 1 0 20332 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 0
transform -1 0 19872 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 0
transform -1 0 18308 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _0945_
timestamp 0
transform 1 0 17020 0 1 18496
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _0946_
timestamp 0
transform 1 0 12972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 0
transform -1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0948_
timestamp 0
transform 1 0 9292 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 0
transform 1 0 9752 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0951_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 0
transform 1 0 21160 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 0
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 0
transform 1 0 9292 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0957_
timestamp 0
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0958_
timestamp 0
transform 1 0 21804 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 0
transform -1 0 21712 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 0
transform 1 0 21988 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 0
transform -1 0 21712 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _0962_
timestamp 0
transform 1 0 14352 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0963_
timestamp 0
transform 1 0 11960 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0964_
timestamp 0
transform 1 0 9384 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0965_
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0966_
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0967_
timestamp 0
transform 1 0 9200 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0968_
timestamp 0
transform 1 0 23828 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0969_
timestamp 0
transform -1 0 25852 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 0
transform 1 0 21252 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 0
transform 1 0 25852 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0972_
timestamp 0
transform 1 0 26036 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 0
transform 1 0 25024 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0974_
timestamp 0
transform 1 0 16836 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0975_
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0976_
timestamp 0
transform 1 0 17296 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0977_
timestamp 0
transform -1 0 15180 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0978_
timestamp 0
transform 1 0 12144 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0979_
timestamp 0
transform 1 0 12144 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0980_
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0981_
timestamp 0
transform 1 0 11592 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0982_
timestamp 0
transform 1 0 27416 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0983_
timestamp 0
transform 1 0 27324 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 0
transform 1 0 15732 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 0
transform 1 0 11868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 0
transform -1 0 14168 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 0
transform 1 0 25392 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 0
transform -1 0 27784 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 0
transform 1 0 14168 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 0
transform 1 0 11500 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 0
transform 1 0 9292 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 0
transform 1 0 22908 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 0
transform 1 0 8740 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 0
transform -1 0 26036 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 0
transform 1 0 6900 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 0
transform 1 0 5612 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 0
transform 1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 0
transform 1 0 17940 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 0
transform 1 0 6900 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 0
transform -1 0 20424 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 0
transform 1 0 19228 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 0
transform 1 0 5520 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 0
transform 1 0 4784 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 0
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 0
transform 1 0 5060 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 0
transform 1 0 20424 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 0
transform 1 0 20056 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 0
transform 1 0 20056 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 0
transform 1 0 5428 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 0
transform 1 0 5060 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 0
transform 1 0 19412 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 0
transform 1 0 5428 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 0
transform -1 0 16560 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 0
transform 1 0 12512 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 0
transform 1 0 11868 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 0
transform 1 0 12880 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 0
transform 1 0 12236 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 0
transform -1 0 26220 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 0
transform -1 0 25944 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 0
transform 1 0 12420 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 0
transform 1 0 9476 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 0
transform 1 0 9200 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 0
transform 1 0 22172 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 0
transform 1 0 8740 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 0
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 0
transform 1 0 9936 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 0
transform 1 0 8004 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 0
transform 1 0 8188 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 0
transform 1 0 23276 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 0
transform 1 0 7912 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 0
transform -1 0 26036 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 0
transform 1 0 24288 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 0
transform 1 0 14628 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 0
transform -1 0 15732 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 0
transform 1 0 11684 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 0
transform 1 0 12052 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 0
transform 1 0 17388 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 0
transform 1 0 13064 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 0
transform 1 0 17480 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 0
transform 1 0 17480 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 0
transform -1 0 16192 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 0
transform 1 0 9568 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 0
transform 1 0 9568 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 0
transform 1 0 17296 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 0
transform 1 0 10672 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 0
transform 1 0 17204 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 0
transform 1 0 17020 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 0
transform 1 0 2024 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 0
transform 1 0 3312 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 0
transform 1 0 2392 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 0
transform 1 0 1932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 0
transform 1 0 14904 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 0
transform 1 0 2208 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 0
transform 1 0 16192 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 0
transform 1 0 1932 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 0
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 0
transform 1 0 1932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 0
transform 1 0 14720 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 0
transform 1 0 2116 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 0
transform 1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 0
transform -1 0 13616 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 0
transform 1 0 7360 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 0
transform 1 0 6992 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 0
transform 1 0 7820 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 0
transform 1 0 21712 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 0
transform 1 0 7360 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 0
transform -1 0 25852 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 0
transform 1 0 22632 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 0
transform 1 0 5704 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 0
transform 1 0 3864 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 0
transform 1 0 3680 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 0
transform 1 0 20240 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 0
transform 1 0 3864 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 0
transform 1 0 20240 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 0
transform 1 0 19872 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 0
transform 1 0 12420 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 0
transform 1 0 8280 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 0
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 0
transform 1 0 20700 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 0
transform 1 0 8740 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 0
transform 1 0 21712 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 16560 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk
timestamp 0
transform -1 0 9292 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 0
transform 1 0 10396 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 0
transform -1 0 8832 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 0
transform 1 0 10396 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 0
transform -1 0 18860 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 0
transform -1 0 21712 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 0
transform -1 0 20240 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 0
transform -1 0 8832 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 0
transform 1 0 10212 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 0
transform -1 0 9016 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 0
transform 1 0 10396 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 0
transform 1 0 17848 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 0
transform 1 0 20424 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 0
transform -1 0 17940 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 0
transform 1 0 19136 0 -1 26112
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_105
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_175
timestamp 0
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_187
timestamp 0
transform 1 0 18308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_195
timestamp 0
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_233
timestamp 0
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_240
timestamp 0
transform 1 0 23184 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_303
timestamp 0
transform 1 0 28980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 0
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_89
timestamp 0
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_114
timestamp 0
transform 1 0 11592 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_152
timestamp 0
transform 1 0 15088 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_158
timestamp 0
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_175
timestamp 0
transform 1 0 17204 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_200
timestamp 0
transform 1 0 19504 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_212
timestamp 0
transform 1 0 20608 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_224
timestamp 0
transform 1 0 21712 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_236
timestamp 0
transform 1 0 22816 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_248
timestamp 0
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_286
timestamp 0
transform 1 0 27416 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_298
timestamp 0
transform 1 0 28520 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_306
timestamp 0
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_156
timestamp 0
transform 1 0 15456 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_179
timestamp 0
transform 1 0 17572 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_196
timestamp 0
transform 1 0 19136 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_208
timestamp 0
transform 1 0 20240 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_220
timestamp 0
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_301
timestamp 0
transform 1 0 28796 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_313
timestamp 0
transform 1 0 29900 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_106
timestamp 0
transform 1 0 10856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_114
timestamp 0
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_157
timestamp 0
transform 1 0 15548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_171
timestamp 0
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_186
timestamp 0
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 0
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_278
timestamp 0
transform 1 0 26680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_297
timestamp 0
transform 1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_305
timestamp 0
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_87
timestamp 0
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_104
timestamp 0
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_121
timestamp 0
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_155
timestamp 0
transform 1 0 15364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_217
timestamp 0
transform 1 0 21068 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 0
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_234
timestamp 0
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_253
timestamp 0
transform 1 0 24380 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_287
timestamp 0
transform 1 0 27508 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_299
timestamp 0
transform 1 0 28612 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_311
timestamp 0
transform 1 0 29716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_323
timestamp 0
transform 1 0 30820 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 0
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 0
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_88
timestamp 0
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_92
timestamp 0
transform 1 0 9568 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_119
timestamp 0
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_131
timestamp 0
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_157
timestamp 0
transform 1 0 15548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_169
timestamp 0
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_181
timestamp 0
transform 1 0 17756 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_190
timestamp 0
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_206
timestamp 0
transform 1 0 20056 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_212
timestamp 0
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 0
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_286
timestamp 0
transform 1 0 27416 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_298
timestamp 0
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 0
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_77
timestamp 0
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_118
timestamp 0
transform 1 0 11960 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_130
timestamp 0
transform 1 0 13064 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_154
timestamp 0
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 0
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_177
timestamp 0
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_276
timestamp 0
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 0
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 0
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_317
timestamp 0
transform 1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_66
timestamp 0
transform 1 0 7176 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 0
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_111
timestamp 0
transform 1 0 11316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_123
timestamp 0
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 0
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_185
timestamp 0
transform 1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_214
timestamp 0
transform 1 0 20792 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_227
timestamp 0
transform 1 0 21988 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_236
timestamp 0
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 0
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_266
timestamp 0
transform 1 0 25576 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_278
timestamp 0
transform 1 0 26680 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_290
timestamp 0
transform 1 0 27784 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_302
timestamp 0
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_321
timestamp 0
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 0
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 0
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 0
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 0
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 0
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 0
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 0
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 0
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 0
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 0
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_317
timestamp 0
transform 1 0 30268 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 0
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_68
timestamp 0
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_129
timestamp 0
transform 1 0 12972 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 0
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_188
timestamp 0
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 0
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 0
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 0
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 0
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 0
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 0
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 0
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_11
timestamp 0
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_46
timestamp 0
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_106
timestamp 0
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_163
timestamp 0
transform 1 0 16100 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_185
timestamp 0
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_196
timestamp 0
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_218
timestamp 0
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_225
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_252
timestamp 0
transform 1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_271
timestamp 0
transform 1 0 26036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 0
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_317
timestamp 0
transform 1 0 30268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 0
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_40
timestamp 0
transform 1 0 4784 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_46
timestamp 0
transform 1 0 5336 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 0
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_180
timestamp 0
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_275
timestamp 0
transform 1 0 26404 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_287
timestamp 0
transform 1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_299
timestamp 0
transform 1 0 28612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_321
timestamp 0
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 0
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_76
timestamp 0
transform 1 0 8096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_98
timestamp 0
transform 1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_126
timestamp 0
transform 1 0 12696 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_138
timestamp 0
transform 1 0 13800 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_150
timestamp 0
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_158
timestamp 0
transform 1 0 15640 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 0
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_179
timestamp 0
transform 1 0 17572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 0
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_244
timestamp 0
transform 1 0 23552 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_276
timestamp 0
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 0
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 0
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_317
timestamp 0
transform 1 0 30268 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_38
timestamp 0
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_47
timestamp 0
transform 1 0 5428 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_59
timestamp 0
transform 1 0 6532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_74
timestamp 0
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 0
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 0
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_103
timestamp 0
transform 1 0 10580 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_115
timestamp 0
transform 1 0 11684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_127
timestamp 0
transform 1 0 12788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_185
timestamp 0
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 0
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_216
timestamp 0
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_228
timestamp 0
transform 1 0 22080 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_236
timestamp 0
transform 1 0 22816 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_244
timestamp 0
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_272
timestamp 0
transform 1 0 26128 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_284
timestamp 0
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_296
timestamp 0
transform 1 0 28336 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 0
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_321
timestamp 0
transform 1 0 30636 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_19
timestamp 0
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_23
timestamp 0
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 0
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_103
timestamp 0
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 0
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 0
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 0
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_249
timestamp 0
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_258
timestamp 0
transform 1 0 24840 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_270
timestamp 0
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 0
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 0
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_317
timestamp 0
transform 1 0 30268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_11
timestamp 0
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_39
timestamp 0
transform 1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_50
timestamp 0
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_62
timestamp 0
transform 1 0 6808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_74
timestamp 0
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_118
timestamp 0
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_144
timestamp 0
transform 1 0 14352 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_156
timestamp 0
transform 1 0 15456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_160
timestamp 0
transform 1 0 15824 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_208
timestamp 0
transform 1 0 20240 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_220
timestamp 0
transform 1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_224
timestamp 0
transform 1 0 21712 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_234
timestamp 0
transform 1 0 22632 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_246
timestamp 0
transform 1 0 23736 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_277
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_285
timestamp 0
transform 1 0 27324 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_297
timestamp 0
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 0
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 0
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_321
timestamp 0
transform 1 0 30636 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_9
timestamp 0
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_21
timestamp 0
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_32
timestamp 0
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_44
timestamp 0
transform 1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_117
timestamp 0
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_159
timestamp 0
transform 1 0 15732 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_192
timestamp 0
transform 1 0 18768 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_210
timestamp 0
transform 1 0 20424 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_218
timestamp 0
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_244
timestamp 0
transform 1 0 23552 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_256
timestamp 0
transform 1 0 24656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 0
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_317
timestamp 0
transform 1 0 30268 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_76
timestamp 0
transform 1 0 8096 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_80
timestamp 0
transform 1 0 8464 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_101
timestamp 0
transform 1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_116
timestamp 0
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_126
timestamp 0
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_186
timestamp 0
transform 1 0 18216 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_219
timestamp 0
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_269
timestamp 0
transform 1 0 25852 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_281
timestamp 0
transform 1 0 26956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 0
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_321
timestamp 0
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_25
timestamp 0
transform 1 0 3404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_34
timestamp 0
transform 1 0 4232 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_66
timestamp 0
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_72
timestamp 0
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_84
timestamp 0
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_95
timestamp 0
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_129
timestamp 0
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_138
timestamp 0
transform 1 0 13800 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_150
timestamp 0
transform 1 0 14904 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_162
timestamp 0
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_178
timestamp 0
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_187
timestamp 0
transform 1 0 18308 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_285
timestamp 0
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_294
timestamp 0
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_300
timestamp 0
transform 1 0 28704 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_312
timestamp 0
transform 1 0 29808 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_324
timestamp 0
transform 1 0 30912 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_25
timestamp 0
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_49
timestamp 0
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_67
timestamp 0
transform 1 0 7268 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_94
timestamp 0
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_111
timestamp 0
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_123
timestamp 0
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp 0
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_158
timestamp 0
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_170
timestamp 0
transform 1 0 16744 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_182
timestamp 0
transform 1 0 17848 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 0
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 0
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_270
timestamp 0
transform 1 0 25944 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_282
timestamp 0
transform 1 0 27048 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_294
timestamp 0
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_306
timestamp 0
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_317
timestamp 0
transform 1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 0
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_33
timestamp 0
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 0
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_86
timestamp 0
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 0
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 0
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_124
timestamp 0
transform 1 0 12512 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_136
timestamp 0
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_140
timestamp 0
transform 1 0 13984 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_184
timestamp 0
transform 1 0 18032 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_196
timestamp 0
transform 1 0 19136 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_208
timestamp 0
transform 1 0 20240 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_220
timestamp 0
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_258
timestamp 0
transform 1 0 24840 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_270
timestamp 0
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 0
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 0
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_317
timestamp 0
transform 1 0 30268 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_113
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_158
timestamp 0
transform 1 0 15640 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_170
timestamp 0
transform 1 0 16744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_192
timestamp 0
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_273
timestamp 0
transform 1 0 26220 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_290
timestamp 0
transform 1 0 27784 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_302
timestamp 0
transform 1 0 28888 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 0
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_82
timestamp 0
transform 1 0 8648 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_90
timestamp 0
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_95
timestamp 0
transform 1 0 9844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 0
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_144
timestamp 0
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_177
timestamp 0
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_187
timestamp 0
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_196
timestamp 0
transform 1 0 19136 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_208
timestamp 0
transform 1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 0
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_228
timestamp 0
transform 1 0 22080 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_240
timestamp 0
transform 1 0 23184 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_252
timestamp 0
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_264
timestamp 0
transform 1 0 25392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_284
timestamp 0
transform 1 0 27232 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_309
timestamp 0
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_321
timestamp 0
transform 1 0 30636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 0
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 0
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 0
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 0
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_149
timestamp 0
transform 1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_162
timestamp 0
transform 1 0 16008 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_174
timestamp 0
transform 1 0 17112 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 0
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_202
timestamp 0
transform 1 0 19688 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_214
timestamp 0
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_239
timestamp 0
transform 1 0 23092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 0
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_49
timestamp 0
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_74
timestamp 0
transform 1 0 7912 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_108
timestamp 0
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_117
timestamp 0
transform 1 0 11868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_121
timestamp 0
transform 1 0 12236 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_133
timestamp 0
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_145
timestamp 0
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_157
timestamp 0
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 0
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_210
timestamp 0
transform 1 0 20424 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_214
timestamp 0
transform 1 0 20792 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_237
timestamp 0
transform 1 0 22908 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_257
timestamp 0
transform 1 0 24748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_269
timestamp 0
transform 1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_317
timestamp 0
transform 1 0 30268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_11
timestamp 0
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_25
timestamp 0
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_37
timestamp 0
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_49
timestamp 0
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_61
timestamp 0
transform 1 0 6716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_73
timestamp 0
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 0
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_90
timestamp 0
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_118
timestamp 0
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 0
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 0
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_148
timestamp 0
transform 1 0 14720 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_179
timestamp 0
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_187
timestamp 0
transform 1 0 18308 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_205
timestamp 0
transform 1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_216
timestamp 0
transform 1 0 20976 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_228
timestamp 0
transform 1 0 22080 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_234
timestamp 0
transform 1 0 22632 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_260
timestamp 0
transform 1 0 25024 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_268
timestamp 0
transform 1 0 25760 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_47
timestamp 0
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 0
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_82
timestamp 0
transform 1 0 8648 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 0
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_118
timestamp 0
transform 1 0 11960 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_126
timestamp 0
transform 1 0 12696 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_146
timestamp 0
transform 1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_190
timestamp 0
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_201
timestamp 0
transform 1 0 19596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_213
timestamp 0
transform 1 0 20700 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_221
timestamp 0
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_234
timestamp 0
transform 1 0 22632 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_266
timestamp 0
transform 1 0 25576 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 0
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_284
timestamp 0
transform 1 0 27232 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_296
timestamp 0
transform 1 0 28336 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_308
timestamp 0
transform 1 0 29440 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_320
timestamp 0
transform 1 0 30544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_324
timestamp 0
transform 1 0 30912 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_18
timestamp 0
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 0
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 0
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_98
timestamp 0
transform 1 0 10120 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_116
timestamp 0
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_150
timestamp 0
transform 1 0 14904 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_213
timestamp 0
transform 1 0 20700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_238
timestamp 0
transform 1 0 23000 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 0
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_268
timestamp 0
transform 1 0 25760 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_291
timestamp 0
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_303
timestamp 0
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_321
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_7
timestamp 0
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_43
timestamp 0
transform 1 0 5060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_80
timestamp 0
transform 1 0 8464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_107
timestamp 0
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_121
timestamp 0
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_139
timestamp 0
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_187
timestamp 0
transform 1 0 18308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_195
timestamp 0
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_200
timestamp 0
transform 1 0 19504 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_212
timestamp 0
transform 1 0 20608 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_218
timestamp 0
transform 1 0 21160 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_222
timestamp 0
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_244
timestamp 0
transform 1 0 23552 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_254
timestamp 0
transform 1 0 24472 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_265
timestamp 0
transform 1 0 25484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_277
timestamp 0
transform 1 0 26588 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_285
timestamp 0
transform 1 0 27324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_297
timestamp 0
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_309
timestamp 0
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_321
timestamp 0
transform 1 0 30636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_11
timestamp 0
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_46
timestamp 0
transform 1 0 5336 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_58
timestamp 0
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_90
timestamp 0
transform 1 0 9384 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_102
timestamp 0
transform 1 0 10488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_114
timestamp 0
transform 1 0 11592 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_129
timestamp 0
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp 0
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_150
timestamp 0
transform 1 0 14904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_158
timestamp 0
transform 1 0 15640 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_187
timestamp 0
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_220
timestamp 0
transform 1 0 21344 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_228
timestamp 0
transform 1 0 22080 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_240
timestamp 0
transform 1 0 23184 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_264
timestamp 0
transform 1 0 25392 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_276
timestamp 0
transform 1 0 26496 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_288
timestamp 0
transform 1 0 27600 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_300
timestamp 0
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_19
timestamp 0
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_37
timestamp 0
transform 1 0 4508 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_49
timestamp 0
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_153
timestamp 0
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_183
timestamp 0
transform 1 0 17940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_195
timestamp 0
transform 1 0 19044 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_208
timestamp 0
transform 1 0 20240 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_255
timestamp 0
transform 1 0 24564 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_317
timestamp 0
transform 1 0 30268 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_47
timestamp 0
transform 1 0 5428 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_51
timestamp 0
transform 1 0 5796 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_63
timestamp 0
transform 1 0 6900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_75
timestamp 0
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_101
timestamp 0
transform 1 0 10396 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_115
timestamp 0
transform 1 0 11684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_128
timestamp 0
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_170
timestamp 0
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_182
timestamp 0
transform 1 0 17848 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_190
timestamp 0
transform 1 0 18584 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_203
timestamp 0
transform 1 0 19780 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_207
timestamp 0
transform 1 0 20148 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_257
timestamp 0
transform 1 0 24748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_269
timestamp 0
transform 1 0 25852 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_275
timestamp 0
transform 1 0 26404 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_279
timestamp 0
transform 1 0 26772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_291
timestamp 0
transform 1 0 27876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_303
timestamp 0
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_36
timestamp 0
transform 1 0 4416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_66
timestamp 0
transform 1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_72
timestamp 0
transform 1 0 7728 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_76
timestamp 0
transform 1 0 8096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 0
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_146
timestamp 0
transform 1 0 14536 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_154
timestamp 0
transform 1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 0
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_192
timestamp 0
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_204
timestamp 0
transform 1 0 19872 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_210
timestamp 0
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_266
timestamp 0
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 0
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_317
timestamp 0
transform 1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_54
timestamp 0
transform 1 0 6072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_80
timestamp 0
transform 1 0 8464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_89
timestamp 0
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_110
timestamp 0
transform 1 0 11224 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_127
timestamp 0
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_149
timestamp 0
transform 1 0 14812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 0
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_204
timestamp 0
transform 1 0 19872 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_232
timestamp 0
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_240
timestamp 0
transform 1 0 23184 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_244
timestamp 0
transform 1 0 23552 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_257
timestamp 0
transform 1 0 24748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_269
timestamp 0
transform 1 0 25852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_281
timestamp 0
transform 1 0 26956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_293
timestamp 0
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 0
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_64
timestamp 0
transform 1 0 6992 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_72
timestamp 0
transform 1 0 7728 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_108
timestamp 0
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_140
timestamp 0
transform 1 0 13984 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_152
timestamp 0
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_188
timestamp 0
transform 1 0 18400 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_200
timestamp 0
transform 1 0 19504 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_212
timestamp 0
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_231
timestamp 0
transform 1 0 22356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_239
timestamp 0
transform 1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_256
timestamp 0
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_268
timestamp 0
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_317
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_82
timestamp 0
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_92
timestamp 0
transform 1 0 9568 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_100
timestamp 0
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_149
timestamp 0
transform 1 0 14812 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_159
timestamp 0
transform 1 0 15732 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_184
timestamp 0
transform 1 0 18032 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_217
timestamp 0
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_229
timestamp 0
transform 1 0 22172 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_241
timestamp 0
transform 1 0 23276 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_249
timestamp 0
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_257
timestamp 0
transform 1 0 24748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_269
timestamp 0
transform 1 0 25852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_281
timestamp 0
transform 1 0 26956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_293
timestamp 0
transform 1 0 28060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_305
timestamp 0
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_49
timestamp 0
transform 1 0 5612 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_76
timestamp 0
transform 1 0 8096 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_88
timestamp 0
transform 1 0 9200 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_100
timestamp 0
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_138
timestamp 0
transform 1 0 13800 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_151
timestamp 0
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_163
timestamp 0
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_245
timestamp 0
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_252
timestamp 0
transform 1 0 24288 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_264
timestamp 0
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_276
timestamp 0
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_317
timestamp 0
transform 1 0 30268 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 0
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_37
timestamp 0
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_113
timestamp 0
transform 1 0 11500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_120
timestamp 0
transform 1 0 12144 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_149
timestamp 0
transform 1 0 14812 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_160
timestamp 0
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_172
timestamp 0
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_184
timestamp 0
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_232
timestamp 0
transform 1 0 22448 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_236
timestamp 0
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_240
timestamp 0
transform 1 0 23184 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_244
timestamp 0
transform 1 0 23552 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_270
timestamp 0
transform 1 0 25944 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_282
timestamp 0
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_294
timestamp 0
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 0
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_35
timestamp 0
transform 1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_100
timestamp 0
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_131
timestamp 0
transform 1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_135
timestamp 0
transform 1 0 13524 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_180
timestamp 0
transform 1 0 17664 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 0
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_248
timestamp 0
transform 1 0 23920 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 0
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_317
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_9
timestamp 0
transform 1 0 1932 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_21
timestamp 0
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 0
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_101
timestamp 0
transform 1 0 10396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_119
timestamp 0
transform 1 0 12052 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_131
timestamp 0
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_167
timestamp 0
transform 1 0 16468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_229
timestamp 0
transform 1 0 22172 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_250
timestamp 0
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_271
timestamp 0
transform 1 0 26036 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_283
timestamp 0
transform 1 0 27140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_295
timestamp 0
transform 1 0 28244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_321
timestamp 0
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_44
timestamp 0
transform 1 0 5152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_50
timestamp 0
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_64
timestamp 0
transform 1 0 6992 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_72
timestamp 0
transform 1 0 7728 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_86
timestamp 0
transform 1 0 9016 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_120
timestamp 0
transform 1 0 12144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_139
timestamp 0
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_143
timestamp 0
transform 1 0 14260 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_152
timestamp 0
transform 1 0 15088 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_164
timestamp 0
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 0
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_233
timestamp 0
transform 1 0 22540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_245
timestamp 0
transform 1 0 23644 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_263
timestamp 0
transform 1 0 25300 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_275
timestamp 0
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_317
timestamp 0
transform 1 0 30268 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_76
timestamp 0
transform 1 0 8096 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_80
timestamp 0
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_116
timestamp 0
transform 1 0 11776 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_135
timestamp 0
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_149
timestamp 0
transform 1 0 14812 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_161
timestamp 0
transform 1 0 15916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_173
timestamp 0
transform 1 0 17020 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_205
timestamp 0
transform 1 0 19964 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_217
timestamp 0
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_229
timestamp 0
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_241
timestamp 0
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_249
timestamp 0
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 0
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 0
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_49
timestamp 0
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 0
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_144
timestamp 0
transform 1 0 14352 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_156
timestamp 0
transform 1 0 15456 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_207
timestamp 0
transform 1 0 20148 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_219
timestamp 0
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_268
timestamp 0
transform 1 0 25760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_116
timestamp 0
transform 1 0 11776 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_128
timestamp 0
transform 1 0 12880 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_149
timestamp 0
transform 1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_157
timestamp 0
transform 1 0 15548 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_168
timestamp 0
transform 1 0 16560 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_183
timestamp 0
transform 1 0 17940 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_226
timestamp 0
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_238
timestamp 0
transform 1 0 23000 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_246
timestamp 0
transform 1 0 23736 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_269
timestamp 0
transform 1 0 25852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_281
timestamp 0
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_293
timestamp 0
transform 1 0 28060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 0
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_135
timestamp 0
transform 1 0 13524 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_147
timestamp 0
transform 1 0 14628 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_151
timestamp 0
transform 1 0 14996 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_201
timestamp 0
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_222
timestamp 0
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_236
timestamp 0
transform 1 0 22816 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_256
timestamp 0
transform 1 0 24656 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_276
timestamp 0
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 0
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_317
timestamp 0
transform 1 0 30268 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_33
timestamp 0
transform 1 0 4140 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_37
timestamp 0
transform 1 0 4508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_49
timestamp 0
transform 1 0 5612 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_71
timestamp 0
transform 1 0 7636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_117
timestamp 0
transform 1 0 11868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 0
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_149
timestamp 0
transform 1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_157
timestamp 0
transform 1 0 15548 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_175
timestamp 0
transform 1 0 17204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_187
timestamp 0
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_243
timestamp 0
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 0
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_280
timestamp 0
transform 1 0 26864 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_292
timestamp 0
transform 1 0 27968 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_304
timestamp 0
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_88
timestamp 0
transform 1 0 9200 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_100
timestamp 0
transform 1 0 10304 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 0
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_121
timestamp 0
transform 1 0 12236 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_129
timestamp 0
transform 1 0 12972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_141
timestamp 0
transform 1 0 14076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_153
timestamp 0
transform 1 0 15180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_165
timestamp 0
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_169
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_194
timestamp 0
transform 1 0 18952 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_206
timestamp 0
transform 1 0 20056 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_218
timestamp 0
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_232
timestamp 0
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_236
timestamp 0
transform 1 0 22816 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_250
timestamp 0
transform 1 0 24104 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_262
timestamp 0
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_274
timestamp 0
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_47
timestamp 0
transform 1 0 5428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 0
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_94
timestamp 0
transform 1 0 9752 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_105
timestamp 0
transform 1 0 10764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_117
timestamp 0
transform 1 0 11868 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_126
timestamp 0
transform 1 0 12696 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_149
timestamp 0
transform 1 0 14812 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_163
timestamp 0
transform 1 0 16100 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_175
timestamp 0
transform 1 0 17204 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 0
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_223
timestamp 0
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_235
timestamp 0
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_247
timestamp 0
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_47
timestamp 0
transform 1 0 5428 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_60
timestamp 0
transform 1 0 6624 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_72
timestamp 0
transform 1 0 7728 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_90
timestamp 0
transform 1 0 9384 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_129
timestamp 0
transform 1 0 12972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_146
timestamp 0
transform 1 0 14536 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_150
timestamp 0
transform 1 0 14904 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_160
timestamp 0
transform 1 0 15824 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_177
timestamp 0
transform 1 0 17388 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_207
timestamp 0
transform 1 0 20148 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_233
timestamp 0
transform 1 0 22540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_245
timestamp 0
transform 1 0 23644 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_276
timestamp 0
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 0
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_89
timestamp 0
transform 1 0 9292 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_105
timestamp 0
transform 1 0 10764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_113
timestamp 0
transform 1 0 11500 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_123
timestamp 0
transform 1 0 12420 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_135
timestamp 0
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_171
timestamp 0
transform 1 0 16836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_183
timestamp 0
transform 1 0 17940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_206
timestamp 0
transform 1 0 20056 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_217
timestamp 0
transform 1 0 21068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_229
timestamp 0
transform 1 0 22172 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_235
timestamp 0
transform 1 0 22724 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_271
timestamp 0
transform 1 0 26036 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_283
timestamp 0
transform 1 0 27140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_295
timestamp 0
transform 1 0 28244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_7
timestamp 0
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_19
timestamp 0
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_31
timestamp 0
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_43
timestamp 0
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_66
timestamp 0
transform 1 0 7176 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_74
timestamp 0
transform 1 0 7912 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_79
timestamp 0
transform 1 0 8372 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_91
timestamp 0
transform 1 0 9476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_103
timestamp 0
transform 1 0 10580 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 0
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_130
timestamp 0
transform 1 0 13064 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_138
timestamp 0
transform 1 0 13800 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 0
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 0
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 0
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_191
timestamp 0
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_203
timestamp 0
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_211
timestamp 0
transform 1 0 20516 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_221
timestamp 0
transform 1 0 21436 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_234
timestamp 0
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_265
timestamp 0
transform 1 0 25484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_277
timestamp 0
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_66
timestamp 0
transform 1 0 7176 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_102
timestamp 0
transform 1 0 10488 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_136
timestamp 0
transform 1 0 13616 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_169
timestamp 0
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_192
timestamp 0
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_205
timestamp 0
transform 1 0 19964 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_240
timestamp 0
transform 1 0 23184 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_269
timestamp 0
transform 1 0 25852 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_281
timestamp 0
transform 1 0 26956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_293
timestamp 0
transform 1 0 28060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_305
timestamp 0
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_63
timestamp 0
transform 1 0 6900 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_72
timestamp 0
transform 1 0 7728 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_84
timestamp 0
transform 1 0 8832 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_96
timestamp 0
transform 1 0 9936 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_104
timestamp 0
transform 1 0 10672 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_110
timestamp 0
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_130
timestamp 0
transform 1 0 13064 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_142
timestamp 0
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_154
timestamp 0
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 0
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_177
timestamp 0
transform 1 0 17388 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_214
timestamp 0
transform 1 0 20792 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_233
timestamp 0
transform 1 0 22540 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_243
timestamp 0
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_258
timestamp 0
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_270
timestamp 0
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_278
timestamp 0
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_7
timestamp 0
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_19
timestamp 0
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_57
timestamp 0
transform 1 0 6348 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 0
transform 1 0 7728 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_113
timestamp 0
transform 1 0 11500 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_126
timestamp 0
transform 1 0 12696 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 0
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_169
timestamp 0
transform 1 0 16652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_221
timestamp 0
transform 1 0 21436 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_225
timestamp 0
transform 1 0 21804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_237
timestamp 0
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_249
timestamp 0
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_259
timestamp 0
transform 1 0 24932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_271
timestamp 0
transform 1 0 26036 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_279
timestamp 0
transform 1 0 26772 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_281
timestamp 0
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_293
timestamp 0
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_305
timestamp 0
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_315
timestamp 0
transform 1 0 30084 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_323
timestamp 0
transform 1 0 30820 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 18400 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 28428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 26956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 29256 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform -1 0 14904 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform 1 0 11960 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 16468 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 18308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 26220 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 19688 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 23552 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 14536 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 10948 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 15088 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 14812 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 16836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 20700 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 11224 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 10764 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 0
transform -1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 0
transform -1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 0
transform -1 0 11776 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 0
transform 1 0 4968 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 0
transform -1 0 6164 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 0
transform -1 0 26312 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 0
transform -1 0 7912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 0
transform -1 0 16192 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 0
transform -1 0 10672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 0
transform -1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 0
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 0
transform -1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 0
transform -1 0 4508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 0
transform -1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 0
transform -1 0 24564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 0
transform -1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 0
transform -1 0 7912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 0
transform -1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 0
transform -1 0 19504 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 0
transform -1 0 14812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 0
transform -1 0 4140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 0
transform -1 0 5336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 0
transform 1 0 15640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 0
transform -1 0 25300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 0
transform -1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 0
transform -1 0 12420 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 0
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 0
transform -1 0 25484 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 0
transform -1 0 11132 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 0
transform -1 0 26496 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 0
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 0
transform -1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 0
transform -1 0 5612 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 0
transform -1 0 6164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 0
transform -1 0 22632 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 0
transform -1 0 25760 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 0
transform -1 0 14812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 0
transform -1 0 13064 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 0
transform -1 0 17756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 0
transform -1 0 21620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 0
transform -1 0 22540 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 0
transform -1 0 20976 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 0
transform -1 0 10580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 0
transform -1 0 10488 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 0
transform -1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 0
transform -1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 0
transform -1 0 10396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 0
transform -1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 0
transform 1 0 6532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 0
transform -1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 0
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 0
transform -1 0 7912 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 0
transform -1 0 20792 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 0
transform -1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 0
transform -1 0 10672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 0
transform -1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 0
transform -1 0 14076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 0
transform 1 0 14260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 0
transform -1 0 19228 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 0
transform -1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 0
transform -1 0 23460 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 0
transform -1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 0
transform -1 0 11960 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 0
transform -1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 0
transform 1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 0
transform -1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 0
transform -1 0 17572 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 0
transform -1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 0
transform -1 0 10120 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 0
transform -1 0 19964 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 0
transform -1 0 4140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 0
transform -1 0 10488 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 0
transform -1 0 23552 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 0
transform -1 0 19136 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 0
transform -1 0 13892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 0
transform -1 0 23644 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 0
transform -1 0 22540 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 0
transform -1 0 16560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 0
transform -1 0 19044 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 0
transform -1 0 15272 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 0
transform -1 0 11316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 0
transform -1 0 13064 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 0
transform 1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 0
transform -1 0 4968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 0
transform -1 0 22540 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 0
transform -1 0 5336 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 0
transform -1 0 22816 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 0
transform -1 0 9844 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 0
transform -1 0 24840 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 0
transform -1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 0
transform 1 0 13064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 0
transform -1 0 25944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 0
transform -1 0 28152 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 0
transform -1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 0
transform -1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 0
transform -1 0 7176 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 0
transform -1 0 25392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 0
transform -1 0 6256 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 0
transform -1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 0
transform -1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 0
transform -1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 0
transform -1 0 8556 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 0
transform -1 0 9568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 0
transform -1 0 29164 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 0
transform -1 0 7728 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 0
transform -1 0 26496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 0
transform -1 0 24288 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 0
transform -1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 0
transform -1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 0
transform -1 0 25760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 0
transform -1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 0
transform -1 0 23368 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 0
transform -1 0 11592 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 0
transform -1 0 7912 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 0
transform -1 0 26128 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 0
transform -1 0 26864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 0
transform -1 0 14996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 0
transform 1 0 28428 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 0
transform 1 0 7176 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 0
transform 1 0 12328 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 0
transform 1 0 29716 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 0
transform -1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 0
transform -1 0 31004 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  max_cap24
timestamp 0
transform -1 0 22540 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap25
timestamp 0
transform -1 0 18308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap26
timestamp 0
transform -1 0 24748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap28
timestamp 0
transform -1 0 24748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  max_cap29
timestamp 0
transform 1 0 23368 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 0
transform -1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 0
transform -1 0 1932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 0
transform -1 0 11408 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 0
transform 1 0 30452 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 0
transform -1 0 18308 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 0
transform -1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 31280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 31280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 31280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 31280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 31280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 31280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 31280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 31280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 31280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 31280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 31280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 31280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 31280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 31280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 31280 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 31280 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 31280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 31280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 31280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 31280 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 31280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 31280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 31280 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 31280 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 31280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 31280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 31280 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 31280 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 31280 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 31280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 31280 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 31280 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 31280 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 31280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 31280 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 31280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 31280 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 31280 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 31280 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 31280 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 31280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 31280 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 31280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 0
transform -1 0 31280 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 0
transform -1 0 31280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 0
transform -1 0 31280 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 0
transform -1 0 31280 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 0
transform -1 0 31280 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 0
transform -1 0 31280 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 0
transform -1 0 31280 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 0
transform -1 0 31280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 0
transform 1 0 6256 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 0
transform 1 0 11408 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 0
transform 1 0 16560 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 0
transform 1 0 21712 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 0
transform 1 0 26864 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire1
timestamp 0
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire23
timestamp 0
transform -1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  wire27
timestamp 0
transform -1 0 15732 0 1 21760
box -38 -48 406 592
<< labels >>
rlabel metal1 s 16192 31552 16192 31552 4 VGND
rlabel metal2 s 16192 32096 16192 32096 4 VPWR
rlabel metal1 s 21988 15130 21988 15130 4 _0000_
rlabel metal1 s 27225 16558 27225 16558 4 _0001_
rlabel metal1 s 27140 18054 27140 18054 4 _0002_
rlabel metal2 s 26634 19550 26634 19550 4 _0003_
rlabel metal2 s 17894 14178 17894 14178 4 _0004_
rlabel metal2 s 20194 21522 20194 21522 4 _0005_
rlabel metal1 s 18722 3543 18722 3543 4 _0006_
rlabel metal1 s 14950 4250 14950 4250 4 _0007_
rlabel metal1 s 14313 3434 14313 3434 4 _0008_
rlabel metal1 s 13945 11050 13945 11050 4 _0009_
rlabel metal1 s 27508 3706 27508 3706 4 _0010_
rlabel metal1 s 13347 14314 13347 14314 4 _0011_
rlabel metal1 s 29171 15062 29171 15062 4 _0012_
rlabel metal1 s 28612 12614 28612 12614 4 _0013_
rlabel metal1 s 14474 13974 14474 13974 4 _0014_
rlabel metal1 s 12093 8534 12093 8534 4 _0015_
rlabel metal1 s 9747 3434 9747 3434 4 _0016_
rlabel metal1 s 10345 11730 10345 11730 4 _0017_
rlabel metal1 s 24594 5610 24594 5610 4 _0018_
rlabel metal2 s 9614 15266 9614 15266 4 _0019_
rlabel metal1 s 23950 12886 23950 12886 4 _0020_
rlabel metal1 s 25632 8942 25632 8942 4 _0021_
rlabel metal1 s 21390 15402 21390 15402 4 _0022_
rlabel metal1 s 25842 16762 25842 16762 4 _0023_
rlabel metal1 s 26036 17578 26036 17578 4 _0024_
rlabel metal2 s 25346 19108 25346 19108 4 _0025_
rlabel metal1 s 17342 14450 17342 14450 4 _0026_
rlabel metal1 s 18124 4114 18124 4114 4 _0027_
rlabel metal1 s 14076 4658 14076 4658 4 _0028_
rlabel metal1 s 12328 4658 12328 4658 4 _0029_
rlabel metal1 s 12098 11798 12098 11798 4 _0030_
rlabel metal1 s 27002 4692 27002 4692 4 _0031_
rlabel metal2 s 12466 14484 12466 14484 4 _0032_
rlabel metal1 s 27554 15538 27554 15538 4 _0033_
rlabel metal1 s 27462 11322 27462 11322 4 _0034_
rlabel metal1 s 16049 3502 16049 3502 4 _0035_
rlabel metal1 s 14014 5610 14014 5610 4 _0036_
rlabel metal2 s 12466 4556 12466 4556 4 _0037_
rlabel metal1 s 13948 11730 13948 11730 4 _0038_
rlabel metal1 s 25514 5270 25514 5270 4 _0039_
rlabel metal2 s 12190 15674 12190 15674 4 _0040_
rlabel metal1 s 27374 14314 27374 14314 4 _0041_
rlabel metal1 s 26900 11730 26900 11730 4 _0042_
rlabel metal1 s 14198 14314 14198 14314 4 _0043_
rlabel metal1 s 11576 7786 11576 7786 4 _0044_
rlabel metal2 s 9609 4114 9609 4114 4 _0045_
rlabel metal1 s 9006 11118 9006 11118 4 _0046_
rlabel metal1 s 23455 5202 23455 5202 4 _0047_
rlabel metal1 s 8862 16150 8862 16150 4 _0048_
rlabel metal1 s 23598 12614 23598 12614 4 _0049_
rlabel metal1 s 25816 8466 25816 8466 4 _0050_
rlabel metal1 s 6746 15402 6746 15402 4 _0051_
rlabel metal1 s 6568 8466 6568 8466 4 _0052_
rlabel metal1 s 5648 5678 5648 5678 4 _0053_
rlabel metal1 s 5239 12818 5239 12818 4 _0054_
rlabel metal1 s 18308 5882 18308 5882 4 _0055_
rlabel metal1 s 6256 17306 6256 17306 4 _0056_
rlabel metal1 s 20204 11730 20204 11730 4 _0057_
rlabel metal1 s 19136 9146 19136 9146 4 _0058_
rlabel metal1 s 6113 28458 6113 28458 4 _0059_
rlabel metal2 s 5382 22882 5382 22882 4 _0060_
rlabel metal2 s 5566 20230 5566 20230 4 _0061_
rlabel metal2 s 5474 25058 5474 25058 4 _0062_
rlabel metal2 s 21390 26520 21390 26520 4 _0063_
rlabel metal1 s 6302 27642 6302 27642 4 _0064_
rlabel metal1 s 20178 27030 20178 27030 4 _0065_
rlabel metal1 s 20787 23766 20787 23766 4 _0066_
rlabel metal2 s 5842 15266 5842 15266 4 _0067_
rlabel metal1 s 6108 8942 6108 8942 4 _0068_
rlabel metal1 s 6568 6290 6568 6290 4 _0069_
rlabel metal2 s 5566 12002 5566 12002 4 _0070_
rlabel metal1 s 19632 6290 19632 6290 4 _0071_
rlabel metal1 s 5837 17578 5837 17578 4 _0072_
rlabel metal1 s 19545 12138 19545 12138 4 _0073_
rlabel metal1 s 20562 8602 20562 8602 4 _0074_
rlabel metal1 s 16529 27030 16529 27030 4 _0075_
rlabel metal1 s 12634 23018 12634 23018 4 _0076_
rlabel metal2 s 12185 20434 12185 20434 4 _0077_
rlabel metal1 s 13105 25942 13105 25942 4 _0078_
rlabel metal1 s 24456 26282 24456 26282 4 _0079_
rlabel metal1 s 12473 27370 12473 27370 4 _0080_
rlabel metal1 s 26097 27030 26097 27030 4 _0081_
rlabel metal1 s 26097 23018 26097 23018 4 _0082_
rlabel metal2 s 12732 18326 12732 18326 4 _0083_
rlabel metal1 s 9598 8874 9598 8874 4 _0084_
rlabel metal1 s 9430 4794 9430 4794 4 _0085_
rlabel metal1 s 9000 12138 9000 12138 4 _0086_
rlabel metal2 s 22310 5338 22310 5338 4 _0087_
rlabel metal2 s 9154 17000 9154 17000 4 _0088_
rlabel metal1 s 21873 12954 21873 12954 4 _0089_
rlabel metal1 s 23225 8466 23225 8466 4 _0090_
rlabel metal1 s 10580 28730 10580 28730 4 _0091_
rlabel metal1 s 8367 23766 8367 23766 4 _0092_
rlabel metal2 s 8505 20434 8505 20434 4 _0093_
rlabel metal1 s 9000 26282 9000 26282 4 _0094_
rlabel metal1 s 23496 30226 23496 30226 4 _0095_
rlabel metal1 s 8275 29206 8275 29206 4 _0096_
rlabel metal2 s 26266 29410 26266 29410 4 _0097_
rlabel metal1 s 24410 23766 24410 23766 4 _0098_
rlabel metal1 s 14904 29274 14904 29274 4 _0099_
rlabel metal2 s 13846 23970 13846 23970 4 _0100_
rlabel metal2 s 12558 21318 12558 21318 4 _0101_
rlabel metal1 s 12328 24922 12328 24922 4 _0102_
rlabel metal1 s 17480 28186 17480 28186 4 _0103_
rlabel metal1 s 13110 28730 13110 28730 4 _0104_
rlabel metal1 s 17797 28050 17797 28050 4 _0105_
rlabel metal2 s 17618 24310 17618 24310 4 _0106_
rlabel metal1 s 14152 30634 14152 30634 4 _0107_
rlabel metal1 s 15972 23698 15972 23698 4 _0108_
rlabel metal1 s 9614 21862 9614 21862 4 _0109_
rlabel metal1 s 9690 25194 9690 25194 4 _0110_
rlabel metal1 s 17280 30634 17280 30634 4 _0111_
rlabel metal2 s 10989 30702 10989 30702 4 _0112_
rlabel metal1 s 17470 30226 17470 30226 4 _0113_
rlabel metal1 s 17337 24174 17337 24174 4 _0114_
rlabel metal1 s 2100 15402 2100 15402 4 _0115_
rlabel metal1 s 3721 10710 3721 10710 4 _0116_
rlabel metal2 s 2714 8262 2714 8262 4 _0117_
rlabel metal1 s 2054 13226 2054 13226 4 _0118_
rlabel metal1 s 14934 7446 14934 7446 4 _0119_
rlabel metal1 s 2571 18666 2571 18666 4 _0120_
rlabel metal1 s 16872 11730 16872 11730 4 _0121_
rlabel metal1 s 16406 8874 16406 8874 4 _0122_
rlabel metal2 s 2346 16286 2346 16286 4 _0123_
rlabel metal2 s 2990 10914 2990 10914 4 _0124_
rlabel metal1 s 2295 8874 2295 8874 4 _0125_
rlabel metal2 s 2249 12818 2249 12818 4 _0126_
rlabel metal2 s 15037 7854 15037 7854 4 _0127_
rlabel metal1 s 2484 17850 2484 17850 4 _0128_
rlabel metal1 s 16130 11050 16130 11050 4 _0129_
rlabel metal1 s 16728 8534 16728 8534 4 _0130_
rlabel metal2 s 12834 30328 12834 30328 4 _0131_
rlabel metal1 s 7820 22746 7820 22746 4 _0132_
rlabel metal2 s 7498 20706 7498 20706 4 _0133_
rlabel metal1 s 8188 25466 8188 25466 4 _0134_
rlabel metal1 s 21932 30702 21932 30702 4 _0135_
rlabel metal2 s 8142 30498 8142 30498 4 _0136_
rlabel metal1 s 24798 30634 24798 30634 4 _0137_
rlabel metal1 s 22908 23290 22908 23290 4 _0138_
rlabel metal1 s 5826 30634 5826 30634 4 _0139_
rlabel metal1 s 4227 22678 4227 22678 4 _0140_
rlabel metal2 s 4186 20706 4186 20706 4 _0141_
rlabel metal2 s 3997 24786 3997 24786 4 _0142_
rlabel metal1 s 20695 29206 20695 29206 4 _0143_
rlabel metal1 s 4462 27642 4462 27642 4 _0144_
rlabel metal2 s 20557 30634 20557 30634 4 _0145_
rlabel metal1 s 20138 24106 20138 24106 4 _0146_
rlabel metal1 s 12374 17544 12374 17544 4 _0147_
rlabel metal2 s 8873 8466 8873 8466 4 _0148_
rlabel metal2 s 8970 6086 8970 6086 4 _0149_
rlabel metal1 s 7953 13226 7953 13226 4 _0150_
rlabel metal2 s 21017 5678 21017 5678 4 _0151_
rlabel metal1 s 9103 18326 9103 18326 4 _0152_
rlabel metal1 s 21712 11866 21712 11866 4 _0153_
rlabel metal1 s 21758 8602 21758 8602 4 _0154_
rlabel metal1 s 18768 16082 18768 16082 4 _0155_
rlabel metal2 s 18722 14960 18722 14960 4 _0156_
rlabel metal1 s 21114 20944 21114 20944 4 _0157_
rlabel metal1 s 23598 17204 23598 17204 4 _0158_
rlabel metal2 s 12100 8942 12100 8942 4 _0159_
rlabel metal2 s 21114 19516 21114 19516 4 _0160_
rlabel metal1 s 21206 18938 21206 18938 4 _0161_
rlabel metal1 s 21022 18802 21022 18802 4 _0162_
rlabel metal1 s 21896 17646 21896 17646 4 _0163_
rlabel metal2 s 20746 16864 20746 16864 4 _0164_
rlabel metal1 s 21114 20502 21114 20502 4 _0165_
rlabel metal1 s 25162 20536 25162 20536 4 _0166_
rlabel metal1 s 14490 16490 14490 16490 4 _0167_
rlabel metal1 s 21114 19754 21114 19754 4 _0168_
rlabel metal3 s 14766 18717 14766 18717 4 _0169_
rlabel metal1 s 14858 18870 14858 18870 4 _0170_
rlabel metal1 s 23644 9554 23644 9554 4 _0171_
rlabel metal1 s 24472 9690 24472 9690 4 _0172_
rlabel metal2 s 22024 16966 22024 16966 4 _0173_
rlabel metal1 s 21988 20434 21988 20434 4 _0174_
rlabel metal2 s 21208 12818 21208 12818 4 _0175_
rlabel metal2 s 21390 17850 21390 17850 4 _0176_
rlabel metal2 s 21022 8262 21022 8262 4 _0177_
rlabel metal1 s 20792 19414 20792 19414 4 _0178_
rlabel metal1 s 18906 8432 18906 8432 4 _0179_
rlabel metal1 s 18216 20842 18216 20842 4 _0180_
rlabel metal1 s 19090 8432 19090 8432 4 _0181_
rlabel metal1 s 21666 9622 21666 9622 4 _0182_
rlabel metal1 s 23736 21114 23736 21114 4 _0183_
rlabel metal2 s 24242 21420 24242 21420 4 _0184_
rlabel metal2 s 24334 21182 24334 21182 4 _0185_
rlabel metal1 s 23598 23290 23598 23290 4 _0186_
rlabel metal2 s 20562 21692 20562 21692 4 _0187_
rlabel metal1 s 20194 20978 20194 20978 4 _0188_
rlabel metal1 s 21206 23596 21206 23596 4 _0189_
rlabel metal1 s 16560 20910 16560 20910 4 _0190_
rlabel metal2 s 18446 17816 18446 17816 4 _0191_
rlabel metal2 s 23782 23120 23782 23120 4 _0192_
rlabel metal1 s 16008 18326 16008 18326 4 _0193_
rlabel metal1 s 22264 21114 22264 21114 4 _0194_
rlabel metal1 s 21850 21556 21850 21556 4 _0195_
rlabel metal1 s 22540 23290 22540 23290 4 _0196_
rlabel metal2 s 22954 22950 22954 22950 4 _0197_
rlabel metal1 s 25300 10778 25300 10778 4 _0198_
rlabel metal1 s 14168 15878 14168 15878 4 _0199_
rlabel metal1 s 20332 16490 20332 16490 4 _0200_
rlabel metal1 s 17710 16014 17710 16014 4 _0201_
rlabel metal1 s 26818 11118 26818 11118 4 _0202_
rlabel metal1 s 23552 12206 23552 12206 4 _0203_
rlabel metal1 s 24380 13838 24380 13838 4 _0204_
rlabel metal1 s 20562 12818 20562 12818 4 _0205_
rlabel metal2 s 21390 13328 21390 13328 4 _0206_
rlabel metal1 s 23966 28050 23966 28050 4 _0207_
rlabel metal2 s 21942 28849 21942 28849 4 _0208_
rlabel metal1 s 23966 27098 23966 27098 4 _0209_
rlabel metal1 s 23598 28152 23598 28152 4 _0210_
rlabel metal3 s 24495 15164 24495 15164 4 _0211_
rlabel metal1 s 25162 14042 25162 14042 4 _0212_
rlabel metal1 s 25852 15130 25852 15130 4 _0213_
rlabel metal1 s 10488 16558 10488 16558 4 _0214_
rlabel metal2 s 11178 16932 11178 16932 4 _0215_
rlabel metal1 s 7958 17102 7958 17102 4 _0216_
rlabel metal1 s 10074 16966 10074 16966 4 _0217_
rlabel metal1 s 10902 28050 10902 28050 4 _0218_
rlabel metal1 s 10994 27880 10994 27880 4 _0219_
rlabel metal1 s 11684 27982 11684 27982 4 _0220_
rlabel metal1 s 8372 27574 8372 27574 4 _0221_
rlabel metal2 s 11454 19652 11454 19652 4 _0222_
rlabel metal2 s 12282 15470 12282 15470 4 _0223_
rlabel metal1 s 12650 13906 12650 13906 4 _0224_
rlabel metal1 s 23598 6766 23598 6766 4 _0225_
rlabel metal1 s 25254 6732 25254 6732 4 _0226_
rlabel metal1 s 18400 6766 18400 6766 4 _0227_
rlabel metal1 s 19090 6868 19090 6868 4 _0228_
rlabel metal1 s 23322 28050 23322 28050 4 _0229_
rlabel metal2 s 20746 28560 20746 28560 4 _0230_
rlabel metal1 s 23552 27098 23552 27098 4 _0231_
rlabel metal1 s 23184 27642 23184 27642 4 _0232_
rlabel metal3 s 24242 8908 24242 8908 4 _0233_
rlabel metal2 s 26266 5610 26266 5610 4 _0234_
rlabel metal1 s 26082 4692 26082 4692 4 _0235_
rlabel metal1 s 11316 13158 11316 13158 4 _0236_
rlabel metal1 s 11454 12308 11454 12308 4 _0237_
rlabel metal1 s 4462 12954 4462 12954 4 _0238_
rlabel metal1 s 11454 12648 11454 12648 4 _0239_
rlabel metal2 s 11730 25194 11730 25194 4 _0240_
rlabel metal1 s 12052 24378 12052 24378 4 _0241_
rlabel metal2 s 13386 24480 13386 24480 4 _0242_
rlabel metal1 s 11914 24174 11914 24174 4 _0243_
rlabel metal1 s 11730 12206 11730 12206 4 _0244_
rlabel metal1 s 12466 12240 12466 12240 4 _0245_
rlabel metal2 s 15410 12036 15410 12036 4 _0246_
rlabel metal2 s 11362 6154 11362 6154 4 _0247_
rlabel metal1 s 11822 5882 11822 5882 4 _0248_
rlabel metal1 s 7544 6766 7544 6766 4 _0249_
rlabel metal1 s 11132 6086 11132 6086 4 _0250_
rlabel metal1 s 11270 19822 11270 19822 4 _0251_
rlabel metal2 s 11454 20400 11454 20400 4 _0252_
rlabel metal1 s 11868 19890 11868 19890 4 _0253_
rlabel metal1 s 9752 19754 9752 19754 4 _0254_
rlabel metal1 s 11822 19686 11822 19686 4 _0255_
rlabel metal2 s 11914 5338 11914 5338 4 _0256_
rlabel metal1 s 12466 4624 12466 4624 4 _0257_
rlabel metal1 s 11592 8942 11592 8942 4 _0258_
rlabel metal1 s 12328 9146 12328 9146 4 _0259_
rlabel metal1 s 6900 9554 6900 9554 4 _0260_
rlabel metal1 s 12282 9384 12282 9384 4 _0261_
rlabel metal1 s 11910 23086 11910 23086 4 _0262_
rlabel metal1 s 14398 22712 14398 22712 4 _0263_
rlabel metal2 s 12466 23324 12466 23324 4 _0264_
rlabel metal1 s 9706 22474 9706 22474 4 _0265_
rlabel metal2 s 11868 21284 11868 21284 4 _0266_
rlabel metal1 s 12926 5304 12926 5304 4 _0267_
rlabel metal1 s 12742 5134 12742 5134 4 _0268_
rlabel metal1 s 15318 14994 15318 14994 4 _0269_
rlabel metal1 s 16146 14926 16146 14926 4 _0270_
rlabel metal1 s 7958 15028 7958 15028 4 _0271_
rlabel metal1 s 12650 14926 12650 14926 4 _0272_
rlabel metal1 s 15870 28594 15870 28594 4 _0273_
rlabel metal1 s 15548 28730 15548 28730 4 _0274_
rlabel metal1 s 16100 27642 16100 27642 4 _0275_
rlabel metal2 s 15594 28322 15594 28322 4 _0276_
rlabel metal1 s 15778 15606 15778 15606 4 _0277_
rlabel metal2 s 15824 13804 15824 13804 4 _0278_
rlabel metal1 s 17066 4624 17066 4624 4 _0279_
rlabel metal1 s 20102 15334 20102 15334 4 _0280_
rlabel metal1 s 18262 15538 18262 15538 4 _0281_
rlabel metal1 s 17894 14994 17894 14994 4 _0282_
rlabel metal1 s 23046 17578 23046 17578 4 _0283_
rlabel metal2 s 19642 19333 19642 19333 4 _0284_
rlabel metal1 s 18860 14994 18860 14994 4 _0285_
rlabel metal1 s 20470 17644 20470 17644 4 _0286_
rlabel metal1 s 20562 17306 20562 17306 4 _0287_
rlabel metal2 s 20102 17850 20102 17850 4 _0288_
rlabel metal1 s 23506 17748 23506 17748 4 _0289_
rlabel metal1 s 18722 17850 18722 17850 4 _0290_
rlabel metal1 s 18262 20910 18262 20910 4 _0291_
rlabel metal1 s 18492 17170 18492 17170 4 _0292_
rlabel metal1 s 21114 16014 21114 16014 4 _0293_
rlabel metal1 s 24564 17850 24564 17850 4 _0294_
rlabel metal1 s 23506 16660 23506 16660 4 _0295_
rlabel metal1 s 24380 16082 24380 16082 4 _0296_
rlabel metal2 s 23230 16541 23230 16541 4 _0297_
rlabel metal1 s 24794 16218 24794 16218 4 _0298_
rlabel metal1 s 25392 17306 25392 17306 4 _0299_
rlabel metal1 s 23828 16762 23828 16762 4 _0300_
rlabel metal1 s 25346 17204 25346 17204 4 _0301_
rlabel metal1 s 19366 16694 19366 16694 4 _0302_
rlabel metal2 s 21390 16354 21390 16354 4 _0303_
rlabel metal1 s 20976 15470 20976 15470 4 _0304_
rlabel metal1 s 16422 4624 16422 4624 4 _0305_
rlabel metal1 s 14168 13362 14168 13362 4 _0306_
rlabel metal1 s 14490 13498 14490 13498 4 _0307_
rlabel metal2 s 13846 7446 13846 7446 4 _0308_
rlabel metal1 s 11776 8466 11776 8466 4 _0309_
rlabel metal1 s 13754 20366 13754 20366 4 _0310_
rlabel metal1 s 9246 4624 9246 4624 4 _0311_
rlabel metal2 s 12742 11560 12742 11560 4 _0312_
rlabel metal1 s 11270 11322 11270 11322 4 _0313_
rlabel metal2 s 19734 6086 19734 6086 4 _0314_
rlabel metal1 s 24104 5678 24104 5678 4 _0315_
rlabel metal2 s 13202 15402 13202 15402 4 _0316_
rlabel metal1 s 10258 14994 10258 14994 4 _0317_
rlabel metal1 s 20148 27438 20148 27438 4 _0318_
rlabel metal1 s 24012 12818 24012 12818 4 _0319_
rlabel metal1 s 19780 9894 19780 9894 4 _0320_
rlabel metal1 s 26036 8942 26036 8942 4 _0321_
rlabel metal1 s 17802 13872 17802 13872 4 _0322_
rlabel metal2 s 17802 20332 17802 20332 4 _0323_
rlabel metal1 s 17342 20502 17342 20502 4 _0324_
rlabel metal1 s 17526 16592 17526 16592 4 _0325_
rlabel metal1 s 17526 16694 17526 16694 4 _0326_
rlabel metal1 s 15916 4590 15916 4590 4 _0327_
rlabel metal1 s 13616 6290 13616 6290 4 _0328_
rlabel metal1 s 12880 4794 12880 4794 4 _0329_
rlabel metal1 s 15686 11764 15686 11764 4 _0330_
rlabel metal1 s 25254 5202 25254 5202 4 _0331_
rlabel metal1 s 12742 15130 12742 15130 4 _0332_
rlabel metal1 s 26910 14994 26910 14994 4 _0333_
rlabel metal1 s 25944 11730 25944 11730 4 _0334_
rlabel metal1 s 16514 18190 16514 18190 4 _0335_
rlabel metal1 s 16698 16660 16698 16660 4 _0336_
rlabel metal1 s 14260 8398 14260 8398 4 _0337_
rlabel metal2 s 13754 14586 13754 14586 4 _0338_
rlabel metal1 s 12926 8296 12926 8296 4 _0339_
rlabel metal1 s 10028 4590 10028 4590 4 _0340_
rlabel metal1 s 8740 11730 8740 11730 4 _0341_
rlabel metal1 s 23874 5712 23874 5712 4 _0342_
rlabel metal1 s 9384 16082 9384 16082 4 _0343_
rlabel metal1 s 23322 12750 23322 12750 4 _0344_
rlabel metal1 s 26358 8976 26358 8976 4 _0345_
rlabel metal2 s 17710 20128 17710 20128 4 _0346_
rlabel metal1 s 15916 16762 15916 16762 4 _0347_
rlabel metal2 s 20010 7922 20010 7922 4 _0348_
rlabel metal1 s 5198 15572 5198 15572 4 _0349_
rlabel metal1 s 5474 8908 5474 8908 4 _0350_
rlabel metal1 s 5336 6290 5336 6290 4 _0351_
rlabel metal1 s 6394 12920 6394 12920 4 _0352_
rlabel metal1 s 18906 5678 18906 5678 4 _0353_
rlabel metal1 s 6072 17170 6072 17170 4 _0354_
rlabel metal1 s 21206 12240 21206 12240 4 _0355_
rlabel metal1 s 19044 8942 19044 8942 4 _0356_
rlabel metal1 s 15870 18394 15870 18394 4 _0357_
rlabel metal1 s 16468 19822 16468 19822 4 _0358_
rlabel metal2 s 7038 28934 7038 28934 4 _0359_
rlabel metal1 s 5934 22610 5934 22610 4 _0360_
rlabel metal1 s 6072 19822 6072 19822 4 _0361_
rlabel metal1 s 5658 24820 5658 24820 4 _0362_
rlabel metal1 s 22034 27030 22034 27030 4 _0363_
rlabel metal1 s 6072 27438 6072 27438 4 _0364_
rlabel metal1 s 20148 26962 20148 26962 4 _0365_
rlabel metal2 s 21390 24582 21390 24582 4 _0366_
rlabel metal1 s 16054 18734 16054 18734 4 _0367_
rlabel metal1 s 15686 18666 15686 18666 4 _0368_
rlabel metal1 s 6210 14994 6210 14994 4 _0369_
rlabel metal1 s 5796 8942 5796 8942 4 _0370_
rlabel metal1 s 6256 6766 6256 6766 4 _0371_
rlabel metal1 s 6164 11730 6164 11730 4 _0372_
rlabel metal1 s 17710 6324 17710 6324 4 _0373_
rlabel metal1 s 6256 18258 6256 18258 4 _0374_
rlabel metal1 s 20332 12614 20332 12614 4 _0375_
rlabel metal1 s 21114 8398 21114 8398 4 _0376_
rlabel metal1 s 16008 20570 16008 20570 4 _0377_
rlabel metal1 s 13938 20400 13938 20400 4 _0378_
rlabel metal1 s 16606 26554 16606 26554 4 _0379_
rlabel metal2 s 12282 22916 12282 22916 4 _0380_
rlabel metal1 s 13018 20570 13018 20570 4 _0381_
rlabel metal1 s 12788 25874 12788 25874 4 _0382_
rlabel metal1 s 24150 26010 24150 26010 4 _0383_
rlabel metal2 s 12006 27268 12006 27268 4 _0384_
rlabel metal1 s 26404 26962 26404 26962 4 _0385_
rlabel metal1 s 26358 23698 26358 23698 4 _0386_
rlabel metal1 s 15180 18258 15180 18258 4 _0387_
rlabel metal1 s 15410 18190 15410 18190 4 _0388_
rlabel metal2 s 14122 18292 14122 18292 4 _0389_
rlabel metal1 s 9660 8602 9660 8602 4 _0390_
rlabel metal2 s 9706 5066 9706 5066 4 _0391_
rlabel metal1 s 8970 12614 8970 12614 4 _0392_
rlabel metal1 s 21528 5202 21528 5202 4 _0393_
rlabel metal1 s 9476 16558 9476 16558 4 _0394_
rlabel metal2 s 21482 12988 21482 12988 4 _0395_
rlabel metal1 s 24104 8942 24104 8942 4 _0396_
rlabel metal1 s 19090 20026 19090 20026 4 _0397_
rlabel metal1 s 19228 19142 19228 19142 4 _0398_
rlabel metal2 s 19090 20400 19090 20400 4 _0399_
rlabel metal1 s 19458 21114 19458 21114 4 _0400_
rlabel metal1 s 11132 28526 11132 28526 4 _0401_
rlabel metal1 s 9062 23834 9062 23834 4 _0402_
rlabel metal2 s 9706 20740 9706 20740 4 _0403_
rlabel metal1 s 8970 26010 8970 26010 4 _0404_
rlabel metal1 s 23276 29818 23276 29818 4 _0405_
rlabel metal1 s 8740 28730 8740 28730 4 _0406_
rlabel metal1 s 26450 29070 26450 29070 4 _0407_
rlabel metal1 s 24104 23698 24104 23698 4 _0408_
rlabel metal1 s 17337 21998 17337 21998 4 _0409_
rlabel metal1 s 18768 29070 18768 29070 4 _0410_
rlabel metal1 s 14858 29138 14858 29138 4 _0411_
rlabel metal1 s 13800 23698 13800 23698 4 _0412_
rlabel metal1 s 12972 20910 12972 20910 4 _0413_
rlabel metal1 s 12512 24786 12512 24786 4 _0414_
rlabel metal1 s 17434 28050 17434 28050 4 _0415_
rlabel metal1 s 12972 28526 12972 28526 4 _0416_
rlabel metal1 s 17940 29138 17940 29138 4 _0417_
rlabel metal1 s 17894 23698 17894 23698 4 _0418_
rlabel metal1 s 15916 21522 15916 21522 4 _0419_
rlabel metal2 s 14582 30668 14582 30668 4 _0420_
rlabel metal2 s 14030 30532 14030 30532 4 _0421_
rlabel metal1 s 15916 23290 15916 23290 4 _0422_
rlabel metal1 s 9384 21114 9384 21114 4 _0423_
rlabel metal1 s 9476 24922 9476 24922 4 _0424_
rlabel metal1 s 16882 30702 16882 30702 4 _0425_
rlabel metal1 s 11362 31314 11362 31314 4 _0426_
rlabel metal1 s 17066 30804 17066 30804 4 _0427_
rlabel metal1 s 17480 24786 17480 24786 4 _0428_
rlabel metal1 s 16606 19346 16606 19346 4 _0429_
rlabel metal1 s 17020 19278 17020 19278 4 _0430_
rlabel metal1 s 3450 16014 3450 16014 4 _0431_
rlabel metal2 s 4830 11254 4830 11254 4 _0432_
rlabel metal1 s 3404 7854 3404 7854 4 _0433_
rlabel metal1 s 1702 13396 1702 13396 4 _0434_
rlabel metal1 s 14490 7820 14490 7820 4 _0435_
rlabel metal1 s 3588 18938 3588 18938 4 _0436_
rlabel metal1 s 16330 11798 16330 11798 4 _0437_
rlabel metal1 s 16376 9554 16376 9554 4 _0438_
rlabel metal1 s 16652 17850 16652 17850 4 _0439_
rlabel metal1 s 17618 18156 17618 18156 4 _0440_
rlabel metal1 s 2576 16422 2576 16422 4 _0441_
rlabel metal1 s 3496 10234 3496 10234 4 _0442_
rlabel metal1 s 2576 9554 2576 9554 4 _0443_
rlabel metal1 s 3358 13498 3358 13498 4 _0444_
rlabel metal1 s 15272 8466 15272 8466 4 _0445_
rlabel metal2 s 3634 17850 3634 17850 4 _0446_
rlabel metal2 s 16698 12517 16698 12517 4 _0447_
rlabel metal1 s 16468 8466 16468 8466 4 _0448_
rlabel metal1 s 17342 20876 17342 20876 4 _0449_
rlabel metal1 s 9614 30804 9614 30804 4 _0450_
rlabel metal1 s 11270 30226 11270 30226 4 _0451_
rlabel metal1 s 8510 22610 8510 22610 4 _0452_
rlabel metal1 s 7774 21862 7774 21862 4 _0453_
rlabel metal1 s 8418 25296 8418 25296 4 _0454_
rlabel metal1 s 21620 30022 21620 30022 4 _0455_
rlabel metal1 s 8648 30226 8648 30226 4 _0456_
rlabel metal2 s 24242 31110 24242 31110 4 _0457_
rlabel metal2 s 23138 23290 23138 23290 4 _0458_
rlabel metal1 s 17694 21522 17694 21522 4 _0459_
rlabel metal1 s 21160 28594 21160 28594 4 _0460_
rlabel metal1 s 6026 30362 6026 30362 4 _0461_
rlabel metal1 s 4554 23086 4554 23086 4 _0462_
rlabel metal1 s 4370 20468 4370 20468 4 _0463_
rlabel metal1 s 4232 25262 4232 25262 4 _0464_
rlabel metal1 s 20930 28730 20930 28730 4 _0465_
rlabel metal1 s 4922 27438 4922 27438 4 _0466_
rlabel metal1 s 20700 30362 20700 30362 4 _0467_
rlabel metal1 s 19642 24208 19642 24208 4 _0468_
rlabel metal1 s 17802 18734 17802 18734 4 _0469_
rlabel metal1 s 17250 18666 17250 18666 4 _0470_
rlabel metal2 s 12190 17476 12190 17476 4 _0471_
rlabel metal1 s 9154 8976 9154 8976 4 _0472_
rlabel metal1 s 9476 5678 9476 5678 4 _0473_
rlabel metal1 s 8694 12342 8694 12342 4 _0474_
rlabel metal1 s 21160 6766 21160 6766 4 _0475_
rlabel metal2 s 9338 18292 9338 18292 4 _0476_
rlabel metal1 s 21666 11322 21666 11322 4 _0477_
rlabel metal1 s 21758 8466 21758 8466 4 _0478_
rlabel metal2 s 19688 19516 19688 19516 4 _0479_
rlabel metal3 s 16514 17187 16514 17187 4 clk
rlabel metal3 s 15226 17323 15226 17323 4 clknet_0_clk
rlabel metal1 s 2438 8500 2438 8500 4 clknet_4_0_0_clk
rlabel metal1 s 6578 30702 6578 30702 4 clknet_4_10_0_clk
rlabel metal2 s 12558 24004 12558 24004 4 clknet_4_11_0_clk
rlabel metal1 s 19918 24140 19918 24140 4 clknet_4_12_0_clk
rlabel metal1 s 25576 17714 25576 17714 4 clknet_4_13_0_clk
rlabel metal1 s 16790 26894 16790 26894 4 clknet_4_14_0_clk
rlabel metal1 s 20056 26894 20056 26894 4 clknet_4_15_0_clk
rlabel metal1 s 11730 9554 11730 9554 4 clknet_4_1_0_clk
rlabel metal1 s 2024 13294 2024 13294 4 clknet_4_2_0_clk
rlabel metal1 s 9315 12206 9315 12206 4 clknet_4_3_0_clk
rlabel metal1 s 17342 8466 17342 8466 4 clknet_4_4_0_clk
rlabel metal1 s 21758 5780 21758 5780 4 clknet_4_5_0_clk
rlabel metal2 s 16836 14212 16836 14212 4 clknet_4_6_0_clk
rlabel metal1 s 21850 12852 21850 12852 4 clknet_4_7_0_clk
rlabel metal1 s 2208 18258 2208 18258 4 clknet_4_8_0_clk
rlabel metal2 s 12466 19380 12466 19380 4 clknet_4_9_0_clk
rlabel metal3 s 820 29988 820 29988 4 data_in[0]
rlabel metal2 s 28382 959 28382 959 4 data_in[1]
rlabel metal3 s 1050 5508 1050 5508 4 data_in[2]
rlabel metal3 s 0 17688 800 17808 4 data_in[3]
port 7 nsew
rlabel metal1 s 7222 31790 7222 31790 4 data_in[4]
rlabel metal1 s 12328 31790 12328 31790 4 data_in[5]
rlabel metal1 s 29716 31790 29716 31790 4 data_in[6]
rlabel metal1 s 31142 7854 31142 7854 4 data_in[7]
rlabel metal2 s 22586 1520 22586 1520 4 data_out[0]
rlabel metal2 s 46 1554 46 1554 4 data_out[1]
rlabel metal2 s 5198 959 5198 959 4 data_out[2]
rlabel metal3 s 820 11628 820 11628 4 data_out[3]
rlabel metal2 s 30866 1853 30866 1853 4 data_out[4]
rlabel metal2 s 10994 959 10994 959 4 data_out[5]
rlabel metal1 s 30912 19142 30912 19142 4 data_out[6]
rlabel metal1 s 31096 25466 31096 25466 4 data_out[7]
rlabel metal1 s 17986 31994 17986 31994 4 empty
rlabel metal1 s 24242 31994 24242 31994 4 error
rlabel metal2 s 16790 1520 16790 1520 4 full
rlabel metal1 s 1610 30124 1610 30124 4 net1
rlabel metal2 s 1702 25738 1702 25738 4 net10
rlabel metal1 s 14996 30294 14996 30294 4 net100
rlabel metal1 s 10580 17306 10580 17306 4 net101
rlabel metal1 s 9798 23834 9798 23834 4 net102
rlabel metal1 s 13570 4726 13570 4726 4 net103
rlabel metal1 s 6992 12954 6992 12954 4 net104
rlabel metal1 s 17296 9690 17296 9690 4 net105
rlabel metal1 s 13708 15130 13708 15130 4 net106
rlabel metal1 s 6992 17170 6992 17170 4 net107
rlabel metal1 s 19872 28458 19872 28458 4 net108
rlabel metal1 s 15180 15130 15180 15130 4 net109
rlabel metal2 s 17986 15946 17986 15946 4 net11
rlabel metal1 s 9752 12954 9752 12954 4 net110
rlabel metal1 s 11362 15334 11362 15334 4 net111
rlabel metal1 s 13202 5270 13202 5270 4 net112
rlabel metal1 s 14904 4182 14904 4182 4 net113
rlabel metal1 s 18308 9554 18308 9554 4 net114
rlabel metal1 s 7176 12070 7176 12070 4 net115
rlabel metal1 s 22494 30362 22494 30362 4 net116
rlabel metal1 s 19964 8466 19964 8466 4 net117
rlabel metal1 s 10994 11050 10994 11050 4 net118
rlabel metal2 s 7866 8704 7866 8704 4 net119
rlabel metal1 s 21528 2414 21528 2414 4 net12
rlabel metal1 s 6900 20570 6900 20570 4 net120
rlabel metal1 s 21528 28526 21528 28526 4 net121
rlabel metal1 s 16790 4250 16790 4250 4 net122
rlabel metal1 s 11040 8602 11040 8602 4 net123
rlabel metal1 s 9384 28526 9384 28526 4 net124
rlabel metal1 s 19044 31314 19044 31314 4 net125
rlabel metal1 s 3220 13906 3220 13906 4 net126
rlabel metal1 s 9568 30634 9568 30634 4 net127
rlabel metal1 s 22632 9554 22632 9554 4 net128
rlabel metal1 s 18584 12614 18584 12614 4 net129
rlabel metal1 s 1794 2448 1794 2448 4 net13
rlabel metal1 s 13018 8806 13018 8806 4 net130
rlabel metal1 s 22770 13158 22770 13158 4 net131
rlabel metal1 s 21712 27098 21712 27098 4 net132
rlabel metal1 s 15594 13294 15594 13294 4 net133
rlabel metal1 s 18170 31450 18170 31450 4 net134
rlabel metal1 s 14398 6290 14398 6290 4 net135
rlabel metal1 s 10166 5814 10166 5814 4 net136
rlabel metal2 s 11914 30464 11914 30464 4 net137
rlabel metal2 s 14582 17884 14582 17884 4 net138
rlabel metal1 s 4048 16082 4048 16082 4 net139
rlabel metal1 s 9706 2414 9706 2414 4 net14
rlabel metal1 s 21436 30362 21436 30362 4 net140
rlabel metal1 s 4416 13226 4416 13226 4 net141
rlabel metal1 s 21528 27370 21528 27370 4 net142
rlabel metal1 s 9246 13294 9246 13294 4 net143
rlabel metal1 s 24012 30702 24012 30702 4 net144
rlabel metal1 s 26542 5542 26542 5542 4 net145
rlabel metal1 s 13570 12274 13570 12274 4 net146
rlabel metal1 s 25070 13158 25070 13158 4 net147
rlabel metal1 s 26956 12614 26956 12614 4 net148
rlabel metal1 s 4416 10030 4416 10030 4 net149
rlabel metal1 s 1794 11696 1794 11696 4 net15
rlabel metal1 s 7222 25126 7222 25126 4 net150
rlabel metal1 s 6624 22746 6624 22746 4 net151
rlabel metal1 s 24840 9690 24840 9690 4 net152
rlabel metal1 s 5658 28186 5658 28186 4 net153
rlabel metal1 s 6808 27438 6808 27438 4 net154
rlabel metal1 s 10488 26010 10488 26010 4 net155
rlabel metal1 s 11040 16218 11040 16218 4 net156
rlabel metal1 s 7682 28390 7682 28390 4 net157
rlabel metal1 s 8556 21658 8556 21658 4 net158
rlabel metal1 s 27002 11152 27002 11152 4 net159
rlabel metal1 s 29716 2414 29716 2414 4 net16
rlabel metal1 s 6900 30294 6900 30294 4 net160
rlabel metal1 s 25254 6290 25254 6290 4 net161
rlabel metal1 s 23552 8602 23552 8602 4 net162
rlabel metal2 s 11546 5440 11546 5440 4 net163
rlabel metal1 s 9798 10778 9798 10778 4 net164
rlabel metal1 s 24380 6358 24380 6358 4 net165
rlabel metal1 s 19872 6698 19872 6698 4 net166
rlabel metal1 s 22494 5338 22494 5338 4 net167
rlabel metal1 s 10810 3706 10810 3706 4 net168
rlabel metal1 s 6992 16082 6992 16082 4 net169
rlabel metal1 s 12282 2346 12282 2346 4 net17
rlabel metal1 s 25530 9690 25530 9690 4 net170
rlabel metal1 s 25990 12818 25990 12818 4 net171
rlabel metal1 s 14122 8466 14122 8466 4 net172
rlabel metal1 s 16698 21998 16698 21998 4 net173
rlabel metal1 s 29440 15538 29440 15538 4 net18
rlabel metal1 s 29900 12410 29900 12410 4 net19
rlabel metal1 s 19274 2618 19274 2618 4 net2
rlabel metal1 s 18262 17173 18262 17173 4 net20
rlabel metal3 s 24449 31756 24449 31756 4 net21
rlabel metal1 s 18124 2414 18124 2414 4 net22
rlabel metal2 s 14214 19924 14214 19924 4 net23
rlabel metal1 s 22448 23086 22448 23086 4 net24
rlabel metal1 s 12650 19822 12650 19822 4 net25
rlabel metal2 s 16606 27506 16606 27506 4 net26
rlabel metal1 s 15410 21896 15410 21896 4 net27
rlabel metal1 s 23874 23018 23874 23018 4 net28
rlabel metal1 s 20930 17272 20930 17272 4 net29
rlabel metal1 s 7038 22066 7038 22066 4 net3
rlabel metal2 s 18446 4386 18446 4386 4 net30
rlabel metal1 s 17664 3570 17664 3570 4 net31
rlabel metal1 s 27048 4522 27048 4522 4 net32
rlabel metal1 s 27462 4046 27462 4046 4 net33
rlabel metal1 s 28060 15674 28060 15674 4 net34
rlabel metal1 s 27784 15062 27784 15062 4 net35
rlabel metal1 s 13340 3706 13340 3706 4 net36
rlabel metal1 s 12742 3570 12742 3570 4 net37
rlabel metal2 s 14214 12002 14214 12002 4 net38
rlabel metal1 s 12512 11186 12512 11186 4 net39
rlabel metal1 s 3542 18088 3542 18088 4 net4
rlabel metal1 s 15594 23086 15594 23086 4 net40
rlabel metal1 s 17342 12206 17342 12206 4 net41
rlabel metal1 s 12742 14824 12742 14824 4 net42
rlabel metal2 s 11914 14620 11914 14620 4 net43
rlabel metal1 s 25300 29138 25300 29138 4 net44
rlabel metal1 s 18722 24922 18722 24922 4 net45
rlabel metal1 s 7038 6698 7038 6698 4 net46
rlabel metal1 s 22264 11118 22264 11118 4 net47
rlabel metal1 s 13616 17170 13616 17170 4 net48
rlabel metal1 s 9844 17646 9844 17646 4 net49
rlabel metal1 s 13202 31926 13202 31926 4 net5
rlabel metal1 s 14352 23834 14352 23834 4 net50
rlabel metal1 s 13524 24922 13524 24922 4 net51
rlabel metal1 s 15778 29274 15778 29274 4 net52
rlabel metal1 s 19780 12818 19780 12818 4 net53
rlabel metal1 s 10304 20434 10304 20434 4 net54
rlabel metal1 s 9890 26010 9890 26010 4 net55
rlabel metal1 s 21298 24854 21298 24854 4 net56
rlabel metal1 s 7084 9690 7084 9690 4 net57
rlabel metal2 s 9982 25024 9982 25024 4 net58
rlabel metal1 s 5428 10778 5428 10778 4 net59
rlabel metal2 s 12558 31518 12558 31518 4 net6
rlabel metal1 s 5658 21012 5658 21012 4 net60
rlabel metal1 s 25392 27370 25392 27370 4 net61
rlabel metal1 s 6992 18258 6992 18258 4 net62
rlabel metal1 s 15594 8602 15594 8602 4 net63
rlabel metal1 s 10074 6426 10074 6426 4 net64
rlabel metal1 s 4186 8602 4186 8602 4 net65
rlabel metal1 s 13616 27098 13616 27098 4 net66
rlabel metal1 s 13800 26282 13800 26282 4 net67
rlabel metal1 s 3910 18394 3910 18394 4 net68
rlabel metal1 s 13754 22746 13754 22746 4 net69
rlabel metal1 s 17526 12070 17526 12070 4 net7
rlabel metal1 s 23690 23834 23690 23834 4 net70
rlabel metal1 s 13938 20570 13938 20570 4 net71
rlabel metal1 s 6992 14994 6992 14994 4 net72
rlabel metal1 s 18998 25194 18998 25194 4 net73
rlabel metal1 s 18584 29138 18584 29138 4 net74
rlabel metal1 s 13800 28458 13800 28458 4 net75
rlabel metal1 s 3220 9554 3220 9554 4 net76
rlabel metal1 s 4416 18666 4416 18666 4 net77
rlabel metal1 s 16100 26350 16100 26350 4 net78
rlabel metal1 s 24702 24174 24702 24174 4 net79
rlabel metal1 s 18170 9418 18170 9418 4 net8
rlabel metal1 s 17296 12410 17296 12410 4 net80
rlabel metal1 s 11822 29274 11822 29274 4 net81
rlabel metal1 s 3404 16490 3404 16490 4 net82
rlabel metal1 s 24334 29614 24334 29614 4 net83
rlabel metal2 s 9798 21386 9798 21386 4 net84
rlabel metal1 s 25714 23834 25714 23834 4 net85
rlabel metal1 s 26542 15130 26542 15130 4 net86
rlabel metal1 s 6762 5882 6762 5882 4 net87
rlabel metal1 s 4646 25364 4646 25364 4 net88
rlabel metal1 s 5244 23698 5244 23698 4 net89
rlabel metal1 s 1886 20264 1886 20264 4 net9
rlabel metal1 s 21758 6426 21758 6426 4 net90
rlabel metal1 s 24840 25874 24840 25874 4 net91
rlabel metal1 s 13846 21658 13846 21658 4 net92
rlabel metal1 s 12144 31314 12144 31314 4 net93
rlabel metal1 s 16836 7786 16836 7786 4 net94
rlabel metal1 s 20056 5678 20056 5678 4 net95
rlabel metal2 s 21850 23936 21850 23936 4 net96
rlabel metal1 s 20056 9962 20056 9962 4 net97
rlabel metal1 s 9798 9690 9798 9690 4 net98
rlabel metal1 s 9568 23018 9568 23018 4 net99
rlabel metal3 s 820 23868 820 23868 4 pop
rlabel metal1 s 1426 31790 1426 31790 4 push
rlabel metal1 s 31096 13226 31096 13226 4 rst
rlabel metal1 s 17618 4114 17618 4114 4 stack\[0\]\[0\]
rlabel metal1 s 15364 5882 15364 5882 4 stack\[0\]\[1\]
rlabel metal1 s 14720 4590 14720 4590 4 stack\[0\]\[2\]
rlabel metal1 s 13478 11526 13478 11526 4 stack\[0\]\[3\]
rlabel metal1 s 27048 5134 27048 5134 4 stack\[0\]\[4\]
rlabel metal1 s 13478 15674 13478 15674 4 stack\[0\]\[5\]
rlabel metal1 s 26036 14926 26036 14926 4 stack\[0\]\[6\]
rlabel metal1 s 28244 11866 28244 11866 4 stack\[0\]\[7\]
rlabel metal1 s 4830 15946 4830 15946 4 stack\[10\]\[0\]
rlabel metal2 s 4738 10948 4738 10948 4 stack\[10\]\[1\]
rlabel metal1 s 4416 8534 4416 8534 4 stack\[10\]\[2\]
rlabel metal1 s 3680 13430 3680 13430 4 stack\[10\]\[3\]
rlabel metal1 s 16974 7854 16974 7854 4 stack\[10\]\[4\]
rlabel metal1 s 5198 18836 5198 18836 4 stack\[10\]\[5\]
rlabel metal1 s 18124 11866 18124 11866 4 stack\[10\]\[6\]
rlabel metal1 s 18216 8806 18216 8806 4 stack\[10\]\[7\]
rlabel metal2 s 4370 16388 4370 16388 4 stack\[11\]\[0\]
rlabel metal1 s 4554 11220 4554 11220 4 stack\[11\]\[1\]
rlabel metal1 s 4416 9486 4416 9486 4 stack\[11\]\[2\]
rlabel metal1 s 3634 12886 3634 12886 4 stack\[11\]\[3\]
rlabel metal1 s 16974 7990 16974 7990 4 stack\[11\]\[4\]
rlabel metal1 s 4462 18326 4462 18326 4 stack\[11\]\[5\]
rlabel metal1 s 18032 11730 18032 11730 4 stack\[11\]\[6\]
rlabel metal1 s 18538 8534 18538 8534 4 stack\[11\]\[7\]
rlabel metal1 s 12926 30260 12926 30260 4 stack\[12\]\[0\]
rlabel metal1 s 10350 23188 10350 23188 4 stack\[12\]\[1\]
rlabel metal1 s 9522 21386 9522 21386 4 stack\[12\]\[2\]
rlabel metal1 s 10810 26350 10810 26350 4 stack\[12\]\[3\]
rlabel metal1 s 23230 30906 23230 30906 4 stack\[12\]\[4\]
rlabel metal1 s 9568 30702 9568 30702 4 stack\[12\]\[5\]
rlabel metal1 s 24564 30906 24564 30906 4 stack\[12\]\[6\]
rlabel metal1 s 24242 24378 24242 24378 4 stack\[12\]\[7\]
rlabel metal1 s 7866 30566 7866 30566 4 stack\[13\]\[0\]
rlabel metal2 s 6026 23052 6026 23052 4 stack\[13\]\[1\]
rlabel metal1 s 5612 21454 5612 21454 4 stack\[13\]\[2\]
rlabel metal1 s 5750 24650 5750 24650 4 stack\[13\]\[3\]
rlabel metal1 s 21873 29002 21873 29002 4 stack\[13\]\[4\]
rlabel metal1 s 5704 27914 5704 27914 4 stack\[13\]\[5\]
rlabel metal2 s 21666 29308 21666 29308 4 stack\[13\]\[6\]
rlabel metal2 s 21298 24548 21298 24548 4 stack\[13\]\[7\]
rlabel metal2 s 14398 17340 14398 17340 4 stack\[14\]\[0\]
rlabel metal1 s 10994 8908 10994 8908 4 stack\[14\]\[1\]
rlabel metal1 s 10120 6766 10120 6766 4 stack\[14\]\[2\]
rlabel metal2 s 9706 13668 9706 13668 4 stack\[14\]\[3\]
rlabel metal1 s 22264 6222 22264 6222 4 stack\[14\]\[4\]
rlabel metal1 s 10488 18258 10488 18258 4 stack\[14\]\[5\]
rlabel metal1 s 23138 12070 23138 12070 4 stack\[14\]\[6\]
rlabel metal1 s 23276 9146 23276 9146 4 stack\[14\]\[7\]
rlabel metal2 s 15778 14518 15778 14518 4 stack\[15\]\[0\]
rlabel metal1 s 13754 8908 13754 8908 4 stack\[15\]\[1\]
rlabel metal1 s 11638 3570 11638 3570 4 stack\[15\]\[2\]
rlabel metal1 s 11454 11526 11454 11526 4 stack\[15\]\[3\]
rlabel metal1 s 25300 5882 25300 5882 4 stack\[15\]\[4\]
rlabel metal1 s 10626 15368 10626 15368 4 stack\[15\]\[5\]
rlabel metal1 s 25530 12954 25530 12954 4 stack\[15\]\[6\]
rlabel metal1 s 24748 9146 24748 9146 4 stack\[15\]\[7\]
rlabel metal2 s 15576 14994 15576 14994 4 stack\[1\]\[0\]
rlabel metal1 s 12742 8058 12742 8058 4 stack\[1\]\[1\]
rlabel metal2 s 11454 5678 11454 5678 4 stack\[1\]\[2\]
rlabel metal1 s 10534 11322 10534 11322 4 stack\[1\]\[3\]
rlabel metal1 s 24518 6766 24518 6766 4 stack\[1\]\[4\]
rlabel metal1 s 10700 16558 10700 16558 4 stack\[1\]\[5\]
rlabel metal1 s 25116 12410 25116 12410 4 stack\[1\]\[6\]
rlabel metal1 s 23948 9554 23948 9554 4 stack\[1\]\[7\]
rlabel metal1 s 8096 15674 8096 15674 4 stack\[2\]\[0\]
rlabel metal1 s 7682 8602 7682 8602 4 stack\[2\]\[1\]
rlabel metal1 s 7958 5746 7958 5746 4 stack\[2\]\[2\]
rlabel metal2 s 6008 13294 6008 13294 4 stack\[2\]\[3\]
rlabel metal1 s 20424 6086 20424 6086 4 stack\[2\]\[4\]
rlabel metal1 s 7866 17238 7866 17238 4 stack\[2\]\[5\]
rlabel metal1 s 19090 12852 19090 12852 4 stack\[2\]\[6\]
rlabel metal2 s 20838 9554 20838 9554 4 stack\[2\]\[7\]
rlabel metal1 s 8418 28628 8418 28628 4 stack\[3\]\[0\]
rlabel metal1 s 6624 22542 6624 22542 4 stack\[3\]\[1\]
rlabel metal1 s 6532 20978 6532 20978 4 stack\[3\]\[2\]
rlabel metal1 s 7222 25398 7222 25398 4 stack\[3\]\[3\]
rlabel metal1 s 22540 26894 22540 26894 4 stack\[3\]\[4\]
rlabel metal1 s 8096 27914 8096 27914 4 stack\[3\]\[5\]
rlabel metal1 s 22724 27506 22724 27506 4 stack\[3\]\[6\]
rlabel metal1 s 21781 23562 21781 23562 4 stack\[3\]\[7\]
rlabel metal2 s 7774 15164 7774 15164 4 stack\[4\]\[0\]
rlabel metal2 s 7774 9350 7774 9350 4 stack\[4\]\[1\]
rlabel metal1 s 8188 6834 8188 6834 4 stack\[4\]\[2\]
rlabel metal1 s 7222 12342 7222 12342 4 stack\[4\]\[3\]
rlabel metal1 s 20148 6766 20148 6766 4 stack\[4\]\[4\]
rlabel metal1 s 8004 18190 8004 18190 4 stack\[4\]\[5\]
rlabel metal1 s 20884 12750 20884 12750 4 stack\[4\]\[6\]
rlabel metal1 s 20884 9146 20884 9146 4 stack\[4\]\[7\]
rlabel metal1 s 16100 27438 16100 27438 4 stack\[5\]\[0\]
rlabel metal2 s 13938 23460 13938 23460 4 stack\[5\]\[1\]
rlabel metal1 s 13984 20298 13984 20298 4 stack\[5\]\[2\]
rlabel metal1 s 14490 26010 14490 26010 4 stack\[5\]\[3\]
rlabel metal2 s 25806 26758 25806 26758 4 stack\[5\]\[4\]
rlabel metal2 s 13662 27880 13662 27880 4 stack\[5\]\[5\]
rlabel metal1 s 25484 27098 25484 27098 4 stack\[5\]\[6\]
rlabel metal1 s 25438 23290 25438 23290 4 stack\[5\]\[7\]
rlabel metal2 s 14306 17425 14306 17425 4 stack\[6\]\[0\]
rlabel metal1 s 10948 9078 10948 9078 4 stack\[6\]\[1\]
rlabel metal1 s 10994 6222 10994 6222 4 stack\[6\]\[2\]
rlabel metal1 s 10994 13328 10994 13328 4 stack\[6\]\[3\]
rlabel metal1 s 22862 6290 22862 6290 4 stack\[6\]\[4\]
rlabel metal1 s 10580 17646 10580 17646 4 stack\[6\]\[5\]
rlabel metal1 s 23322 12954 23322 12954 4 stack\[6\]\[6\]
rlabel metal1 s 23552 8330 23552 8330 4 stack\[6\]\[7\]
rlabel metal2 s 12374 29070 12374 29070 4 stack\[7\]\[0\]
rlabel metal1 s 10580 24174 10580 24174 4 stack\[7\]\[1\]
rlabel metal1 s 11086 20468 11086 20468 4 stack\[7\]\[2\]
rlabel metal1 s 10902 26486 10902 26486 4 stack\[7\]\[3\]
rlabel metal1 s 23920 30022 23920 30022 4 stack\[7\]\[4\]
rlabel metal1 s 9660 29614 9660 29614 4 stack\[7\]\[5\]
rlabel metal1 s 25208 29206 25208 29206 4 stack\[7\]\[6\]
rlabel metal1 s 25484 23494 25484 23494 4 stack\[7\]\[7\]
rlabel metal1 s 15640 29478 15640 29478 4 stack\[8\]\[0\]
rlabel metal1 s 14628 24378 14628 24378 4 stack\[8\]\[1\]
rlabel metal2 s 13110 21828 13110 21828 4 stack\[8\]\[2\]
rlabel metal1 s 13478 25160 13478 25160 4 stack\[8\]\[3\]
rlabel metal2 s 19826 28934 19826 28934 4 stack\[8\]\[4\]
rlabel metal1 s 13570 29274 13570 29274 4 stack\[8\]\[5\]
rlabel metal2 s 19366 28492 19366 28492 4 stack\[8\]\[6\]
rlabel metal1 s 20010 24752 20010 24752 4 stack\[8\]\[7\]
rlabel metal1 s 15272 30566 15272 30566 4 stack\[9\]\[0\]
rlabel metal1 s 14950 23834 14950 23834 4 stack\[9\]\[1\]
rlabel metal1 s 11316 21318 11316 21318 4 stack\[9\]\[2\]
rlabel metal1 s 11638 25364 11638 25364 4 stack\[9\]\[3\]
rlabel metal1 s 19274 30906 19274 30906 4 stack\[9\]\[4\]
rlabel metal2 s 12926 30192 12926 30192 4 stack\[9\]\[5\]
rlabel metal1 s 18768 30090 18768 30090 4 stack\[9\]\[6\]
rlabel metal1 s 19550 24684 19550 24684 4 stack\[9\]\[7\]
rlabel metal2 s 23874 15878 23874 15878 4 top\[0\]
rlabel metal1 s 26256 18122 26256 18122 4 top\[1\]
rlabel metal1 s 25668 18054 25668 18054 4 top\[2\]
rlabel metal1 s 24978 19414 24978 19414 4 top\[3\]
rlabel metal1 s 18492 14926 18492 14926 4 top\[4\]
flabel metal5 s 1056 30046 31328 30446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 24046 31328 24446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 18046 31328 18446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 12046 31328 12446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6046 31328 6446 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 28908 2128 29308 32144 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 22908 2128 23308 32144 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16908 2128 17308 32144 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 10908 2128 11308 32144 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4908 2128 5308 32144 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 29306 31328 29706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 23306 31328 23706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 17306 31328 17706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11306 31328 11706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5306 31328 5706 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 28168 2128 28568 32144 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 22168 2128 22568 32144 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 16168 2128 16568 32144 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 10168 2128 10568 32144 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4168 2128 4568 32144 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 31652 31288 32452 31408 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 29928 800 30048 0 FreeSans 600 0 0 0 data_in[0]
port 4 nsew
flabel metal2 s 28354 0 28410 800 0 FreeSans 280 90 0 0 data_in[1]
port 5 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 data_in[2]
port 6 nsew
flabel metal3 s 400 17748 400 17748 0 FreeSans 600 0 0 0 data_in[3]
flabel metal2 s 7102 33796 7158 34596 0 FreeSans 280 90 0 0 data_in[4]
port 8 nsew
flabel metal2 s 12254 33796 12310 34596 0 FreeSans 280 90 0 0 data_in[5]
port 9 nsew
flabel metal2 s 29642 33796 29698 34596 0 FreeSans 280 90 0 0 data_in[6]
port 10 nsew
flabel metal3 s 31652 7488 32452 7608 0 FreeSans 600 0 0 0 data_in[7]
port 11 nsew
flabel metal2 s 22558 0 22614 800 0 FreeSans 280 90 0 0 data_out[0]
port 12 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 data_out[1]
port 13 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 data_out[2]
port 14 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 data_out[3]
port 15 nsew
flabel metal3 s 31652 1368 32452 1488 0 FreeSans 600 0 0 0 data_out[4]
port 16 nsew
flabel metal2 s 10966 0 11022 800 0 FreeSans 280 90 0 0 data_out[5]
port 17 nsew
flabel metal3 s 31652 19048 32452 19168 0 FreeSans 600 0 0 0 data_out[6]
port 18 nsew
flabel metal3 s 31652 25168 32452 25288 0 FreeSans 600 0 0 0 data_out[7]
port 19 nsew
flabel metal2 s 18050 33796 18106 34596 0 FreeSans 280 90 0 0 empty
port 20 nsew
flabel metal2 s 23846 33796 23902 34596 0 FreeSans 280 90 0 0 error
port 21 nsew
flabel metal2 s 16762 0 16818 800 0 FreeSans 280 90 0 0 full
port 22 nsew
flabel metal3 s 0 23808 800 23928 0 FreeSans 600 0 0 0 pop
port 23 nsew
flabel metal2 s 1306 33796 1362 34596 0 FreeSans 280 90 0 0 push
port 24 nsew
flabel metal3 s 31652 12928 32452 13048 0 FreeSans 600 0 0 0 rst
port 25 nsew
<< properties >>
string FIXED_BBOX 0 0 32452 34596
<< end >>
