magic
tech sky130A
magscale 1 2
timestamp 1755431338
<< obsli1 >>
rect 1104 2159 31280 32113
<< obsm1 >>
rect 14 2128 31358 32144
<< metal2 >>
rect 1306 33796 1362 34596
rect 7102 33796 7158 34596
rect 12254 33796 12310 34596
rect 18050 33796 18106 34596
rect 23846 33796 23902 34596
rect 29642 33796 29698 34596
rect 18 0 74 800
rect 5170 0 5226 800
rect 10966 0 11022 800
rect 16762 0 16818 800
rect 22558 0 22614 800
rect 28354 0 28410 800
<< obsm2 >>
rect 20 33740 1250 33796
rect 1418 33740 7046 33796
rect 7214 33740 12198 33796
rect 12366 33740 17994 33796
rect 18162 33740 23790 33796
rect 23958 33740 29586 33796
rect 29754 33740 31354 33796
rect 20 856 31354 33740
rect 130 800 5114 856
rect 5282 800 10910 856
rect 11078 800 16706 856
rect 16874 800 22502 856
rect 22670 800 28298 856
rect 28466 800 31354 856
<< metal3 >>
rect 31652 31288 32452 31408
rect 0 29928 800 30048
rect 31652 25168 32452 25288
rect 0 23808 800 23928
rect 31652 19048 32452 19168
rect 0 17688 800 17808
rect 31652 12928 32452 13048
rect 0 11568 800 11688
rect 31652 7488 32452 7608
rect 0 5448 800 5568
rect 31652 1368 32452 1488
<< obsm3 >>
rect 798 31488 31652 32129
rect 798 31208 31572 31488
rect 798 30128 31652 31208
rect 880 29848 31652 30128
rect 798 25368 31652 29848
rect 798 25088 31572 25368
rect 798 24008 31652 25088
rect 880 23728 31652 24008
rect 798 19248 31652 23728
rect 798 18968 31572 19248
rect 798 17888 31652 18968
rect 880 17608 31652 17888
rect 798 13128 31652 17608
rect 798 12848 31572 13128
rect 798 11768 31652 12848
rect 880 11488 31652 11768
rect 798 7688 31652 11488
rect 798 7408 31572 7688
rect 798 5648 31652 7408
rect 880 5368 31652 5648
rect 798 1568 31652 5368
rect 798 1395 31572 1568
<< metal4 >>
rect 4168 2128 4568 32144
rect 4908 2128 5308 32144
rect 10168 2128 10568 32144
rect 10908 2128 11308 32144
rect 16168 2128 16568 32144
rect 16908 2128 17308 32144
rect 22168 2128 22568 32144
rect 22908 2128 23308 32144
rect 28168 2128 28568 32144
rect 28908 2128 29308 32144
<< obsm4 >>
rect 15331 8739 16088 31789
rect 16648 8739 16828 31789
rect 17388 8739 22088 31789
rect 22648 8739 22828 31789
rect 23388 8739 27909 31789
<< metal5 >>
rect 1056 30046 31328 30446
rect 1056 29306 31328 29706
rect 1056 24046 31328 24446
rect 1056 23306 31328 23706
rect 1056 18046 31328 18446
rect 1056 17306 31328 17706
rect 1056 12046 31328 12446
rect 1056 11306 31328 11706
rect 1056 6046 31328 6446
rect 1056 5306 31328 5706
<< labels >>
rlabel metal4 s 4908 2128 5308 32144 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10908 2128 11308 32144 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16908 2128 17308 32144 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 22908 2128 23308 32144 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 28908 2128 29308 32144 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6046 31328 6446 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12046 31328 12446 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18046 31328 18446 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 24046 31328 24446 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 30046 31328 30446 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4168 2128 4568 32144 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10168 2128 10568 32144 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16168 2128 16568 32144 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22168 2128 22568 32144 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 28168 2128 28568 32144 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5306 31328 5706 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11306 31328 11706 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 17306 31328 17706 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 23306 31328 23706 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 29306 31328 29706 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 31652 31288 32452 31408 6 clk
port 3 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 data_in[0]
port 4 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 data_in[1]
port 5 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 data_in[2]
port 6 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 data_in[3]
port 7 nsew signal input
rlabel metal2 s 7102 33796 7158 34596 6 data_in[4]
port 8 nsew signal input
rlabel metal2 s 12254 33796 12310 34596 6 data_in[5]
port 9 nsew signal input
rlabel metal2 s 29642 33796 29698 34596 6 data_in[6]
port 10 nsew signal input
rlabel metal3 s 31652 7488 32452 7608 6 data_in[7]
port 11 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 data_out[0]
port 12 nsew signal output
rlabel metal2 s 18 0 74 800 6 data_out[1]
port 13 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 data_out[2]
port 14 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 data_out[3]
port 15 nsew signal output
rlabel metal3 s 31652 1368 32452 1488 6 data_out[4]
port 16 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 data_out[5]
port 17 nsew signal output
rlabel metal3 s 31652 19048 32452 19168 6 data_out[6]
port 18 nsew signal output
rlabel metal3 s 31652 25168 32452 25288 6 data_out[7]
port 19 nsew signal output
rlabel metal2 s 18050 33796 18106 34596 6 empty
port 20 nsew signal output
rlabel metal2 s 23846 33796 23902 34596 6 error
port 21 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 full
port 22 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 pop
port 23 nsew signal input
rlabel metal2 s 1306 33796 1362 34596 6 push
port 24 nsew signal input
rlabel metal3 s 31652 12928 32452 13048 6 rst
port 25 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32452 34596
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2350892
string GDS_FILE /openlane/designs/lifo/runs/RUN_2025.08.17_11.46.36/results/signoff/lifo.magic.gds
string GDS_START 321388
<< end >>

